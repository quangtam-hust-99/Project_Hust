module mul_signal
(
    input clk ,reset,
    output [15:0] mul_signal_f1,mul_signal_f2
);
wire clk_sample;
chia_tan #(.N(10),.M(399))div_125k(
    .clk(clk),
    .reset(reset),
    .div_clk(clk_sample)
);
reg [15:0] data_f1,data_f2,fsk_mod;
reg [10:0] count;
wire [31:0] temp_f1,temp_f2;
always @(posedge clk_sample or posedge reset)
begin
  if(reset)
  count<=0;
  else 
  count<=count+1;
end
always @*
case(count)
0	:	data_f1=	864	;
1	:	data_f1=	926	;
2	:	data_f1=	128	;
3	:	data_f1=	-790	;
4	:	data_f1=	-974	;
5	:	data_f1=	-255	;
6	:	data_f1=	700	;
7	:	data_f1=	1005	;
8	:	data_f1=	376	;
9	:	data_f1=	-602	;
10	:	data_f1=	-1022	;
11	:	data_f1=	-494	;
12	:	data_f1=	493	;
13	:	data_f1=	1021	;
14	:	data_f1=	601	;
15	:	data_f1=	-377	;
16	:	data_f1=	-1006	;
17	:	data_f1=	-701	;
18	:	data_f1=	254	;
19	:	data_f1=	973	;
20	:	data_f1=	789	;
21	:	data_f1=	-129	;
22	:	data_f1=	-927	;
23	:	data_f1=	-865	;
24	:	data_f1=	0	;
25	:	data_f1=	864	;
26	:	data_f1=	926	;
27	:	data_f1=	128	;
28	:	data_f1=	-790	;
29	:	data_f1=	-974	;
30	:	data_f1=	-255	;
31	:	data_f1=	700	;
32	:	data_f1=	1005	;
33	:	data_f1=	376	;
34	:	data_f1=	-602	;
35	:	data_f1=	-1022	;
36	:	data_f1=	-494	;
37	:	data_f1=	493	;
38	:	data_f1=	1021	;
39	:	data_f1=	601	;
40	:	data_f1=	-377	;
41	:	data_f1=	-1006	;
42	:	data_f1=	-701	;
43	:	data_f1=	254	;
44	:	data_f1=	973	;
45	:	data_f1=	789	;
46	:	data_f1=	-129	;
47	:	data_f1=	-927	;
48	:	data_f1=	-865	;
49	:	data_f1=	0	;
50	:	data_f1=	864	;
51	:	data_f1=	926	;
52	:	data_f1=	128	;
53	:	data_f1=	-790	;
54	:	data_f1=	-974	;
55	:	data_f1=	-255	;
56	:	data_f1=	700	;
57	:	data_f1=	1005	;
58	:	data_f1=	376	;
59	:	data_f1=	-602	;
60	:	data_f1=	-1022	;
61	:	data_f1=	-494	;
62	:	data_f1=	493	;
63	:	data_f1=	1021	;
64	:	data_f1=	601	;
65	:	data_f1=	-377	;
66	:	data_f1=	-1006	;
67	:	data_f1=	-701	;
68	:	data_f1=	254	;
69	:	data_f1=	973	;
70	:	data_f1=	789	;
71	:	data_f1=	-129	;
72	:	data_f1=	-927	;
73	:	data_f1=	-865	;
74	:	data_f1=	0	;
75	:	data_f1=	864	;
76	:	data_f1=	926	;
77	:	data_f1=	128	;
78	:	data_f1=	-790	;
79	:	data_f1=	-974	;
80	:	data_f1=	-255	;
81	:	data_f1=	700	;
82	:	data_f1=	1005	;
83	:	data_f1=	376	;
84	:	data_f1=	-602	;
85	:	data_f1=	-1022	;
86	:	data_f1=	-494	;
87	:	data_f1=	493	;
88	:	data_f1=	1021	;
89	:	data_f1=	601	;
90	:	data_f1=	-377	;
91	:	data_f1=	-1006	;
92	:	data_f1=	-701	;
93	:	data_f1=	254	;
94	:	data_f1=	973	;
95	:	data_f1=	789	;
96	:	data_f1=	-129	;
97	:	data_f1=	-927	;
98	:	data_f1=	-865	;
99	:	data_f1=	-1	;
100	:	data_f1=	864	;
101	:	data_f1=	926	;
102	:	data_f1=	128	;
103	:	data_f1=	-790	;
104	:	data_f1=	-974	;
105	:	data_f1=	-255	;
106	:	data_f1=	700	;
107	:	data_f1=	1005	;
108	:	data_f1=	376	;
109	:	data_f1=	-602	;
110	:	data_f1=	-1022	;
111	:	data_f1=	-494	;
112	:	data_f1=	493	;
113	:	data_f1=	1021	;
114	:	data_f1=	601	;
115	:	data_f1=	-377	;
116	:	data_f1=	-1006	;
117	:	data_f1=	-701	;
118	:	data_f1=	254	;
119	:	data_f1=	973	;
120	:	data_f1=	789	;
121	:	data_f1=	-129	;
122	:	data_f1=	-927	;
123	:	data_f1=	-865	;
124	:	data_f1=	-1	;
125	:	data_f1=	864	;
126	:	data_f1=	926	;
127	:	data_f1=	128	;
128	:	data_f1=	-790	;
129	:	data_f1=	-974	;
130	:	data_f1=	-255	;
131	:	data_f1=	700	;
132	:	data_f1=	1005	;
133	:	data_f1=	376	;
134	:	data_f1=	-602	;
135	:	data_f1=	-1022	;
136	:	data_f1=	-494	;
137	:	data_f1=	493	;
138	:	data_f1=	1021	;
139	:	data_f1=	601	;
140	:	data_f1=	-377	;
141	:	data_f1=	-1006	;
142	:	data_f1=	-701	;
143	:	data_f1=	254	;
144	:	data_f1=	973	;
145	:	data_f1=	789	;
146	:	data_f1=	-129	;
147	:	data_f1=	-927	;
148	:	data_f1=	-865	;
149	:	data_f1=	0	;
150	:	data_f1=	864	;
151	:	data_f1=	926	;
152	:	data_f1=	128	;
153	:	data_f1=	-790	;
154	:	data_f1=	-974	;
155	:	data_f1=	-255	;
156	:	data_f1=	700	;
157	:	data_f1=	1005	;
158	:	data_f1=	376	;
159	:	data_f1=	-602	;
160	:	data_f1=	-1022	;
161	:	data_f1=	-494	;
162	:	data_f1=	493	;
163	:	data_f1=	1021	;
164	:	data_f1=	601	;
165	:	data_f1=	-377	;
166	:	data_f1=	-1006	;
167	:	data_f1=	-701	;
168	:	data_f1=	254	;
169	:	data_f1=	973	;
170	:	data_f1=	789	;
171	:	data_f1=	-129	;
172	:	data_f1=	-927	;
173	:	data_f1=	-865	;
174	:	data_f1=	0	;
175	:	data_f1=	864	;
176	:	data_f1=	926	;
177	:	data_f1=	128	;
178	:	data_f1=	-790	;
179	:	data_f1=	-974	;
180	:	data_f1=	-255	;
181	:	data_f1=	700	;
182	:	data_f1=	1005	;
183	:	data_f1=	376	;
184	:	data_f1=	-602	;
185	:	data_f1=	-1022	;
186	:	data_f1=	-494	;
187	:	data_f1=	493	;
188	:	data_f1=	1021	;
189	:	data_f1=	601	;
190	:	data_f1=	-377	;
191	:	data_f1=	-1006	;
192	:	data_f1=	-701	;
193	:	data_f1=	254	;
194	:	data_f1=	973	;
195	:	data_f1=	789	;
196	:	data_f1=	-129	;
197	:	data_f1=	-927	;
198	:	data_f1=	-865	;
199	:	data_f1=	-1	;
200	:	data_f1=	864	;
201	:	data_f1=	926	;
202	:	data_f1=	128	;
203	:	data_f1=	-790	;
204	:	data_f1=	-974	;
205	:	data_f1=	-255	;
206	:	data_f1=	700	;
207	:	data_f1=	1005	;
208	:	data_f1=	376	;
209	:	data_f1=	-602	;
210	:	data_f1=	-1022	;
211	:	data_f1=	-494	;
212	:	data_f1=	493	;
213	:	data_f1=	1021	;
214	:	data_f1=	601	;
215	:	data_f1=	-377	;
216	:	data_f1=	-1006	;
217	:	data_f1=	-701	;
218	:	data_f1=	254	;
219	:	data_f1=	973	;
220	:	data_f1=	789	;
221	:	data_f1=	-129	;
222	:	data_f1=	-927	;
223	:	data_f1=	-865	;
224	:	data_f1=	-1	;
225	:	data_f1=	864	;
226	:	data_f1=	926	;
227	:	data_f1=	128	;
228	:	data_f1=	-790	;
229	:	data_f1=	-974	;
230	:	data_f1=	-255	;
231	:	data_f1=	700	;
232	:	data_f1=	1005	;
233	:	data_f1=	376	;
234	:	data_f1=	-602	;
235	:	data_f1=	-1022	;
236	:	data_f1=	-494	;
237	:	data_f1=	493	;
238	:	data_f1=	1021	;
239	:	data_f1=	601	;
240	:	data_f1=	-377	;
241	:	data_f1=	-1006	;
242	:	data_f1=	-701	;
243	:	data_f1=	254	;
244	:	data_f1=	973	;
245	:	data_f1=	789	;
246	:	data_f1=	-129	;
247	:	data_f1=	-927	;
248	:	data_f1=	-865	;
249	:	data_f1=	-1	;
250	:	data_f1=	864	;
251	:	data_f1=	926	;
252	:	data_f1=	128	;
253	:	data_f1=	-790	;
254	:	data_f1=	-974	;
255	:	data_f1=	-255	;
256	:	data_f1=	700	;
257	:	data_f1=	1005	;
258	:	data_f1=	376	;
259	:	data_f1=	-602	;
260	:	data_f1=	-1022	;
261	:	data_f1=	-494	;
262	:	data_f1=	493	;
263	:	data_f1=	1021	;
264	:	data_f1=	601	;
265	:	data_f1=	-377	;
266	:	data_f1=	-1006	;
267	:	data_f1=	-701	;
268	:	data_f1=	254	;
269	:	data_f1=	973	;
270	:	data_f1=	789	;
271	:	data_f1=	-129	;
272	:	data_f1=	-927	;
273	:	data_f1=	-865	;
274	:	data_f1=	0	;
275	:	data_f1=	864	;
276	:	data_f1=	926	;
277	:	data_f1=	128	;
278	:	data_f1=	-790	;
279	:	data_f1=	-974	;
280	:	data_f1=	-255	;
281	:	data_f1=	700	;
282	:	data_f1=	1005	;
283	:	data_f1=	376	;
284	:	data_f1=	-602	;
285	:	data_f1=	-1022	;
286	:	data_f1=	-494	;
287	:	data_f1=	493	;
288	:	data_f1=	1021	;
289	:	data_f1=	601	;
290	:	data_f1=	-377	;
291	:	data_f1=	-1006	;
292	:	data_f1=	-701	;
293	:	data_f1=	254	;
294	:	data_f1=	973	;
295	:	data_f1=	789	;
296	:	data_f1=	-129	;
297	:	data_f1=	-927	;
298	:	data_f1=	-865	;
299	:	data_f1=	-1	;
300	:	data_f1=	864	;
301	:	data_f1=	926	;
302	:	data_f1=	128	;
303	:	data_f1=	-790	;
304	:	data_f1=	-974	;
305	:	data_f1=	-255	;
306	:	data_f1=	700	;
307	:	data_f1=	1005	;
308	:	data_f1=	376	;
309	:	data_f1=	-602	;
310	:	data_f1=	-1022	;
311	:	data_f1=	-494	;
312	:	data_f1=	493	;
313	:	data_f1=	1021	;
314	:	data_f1=	601	;
315	:	data_f1=	-377	;
316	:	data_f1=	-1006	;
317	:	data_f1=	-701	;
318	:	data_f1=	254	;
319	:	data_f1=	973	;
320	:	data_f1=	789	;
321	:	data_f1=	-129	;
322	:	data_f1=	-927	;
323	:	data_f1=	-865	;
324	:	data_f1=	0	;
325	:	data_f1=	864	;
326	:	data_f1=	926	;
327	:	data_f1=	128	;
328	:	data_f1=	-790	;
329	:	data_f1=	-974	;
330	:	data_f1=	-255	;
331	:	data_f1=	700	;
332	:	data_f1=	1005	;
333	:	data_f1=	376	;
334	:	data_f1=	-602	;
335	:	data_f1=	-1022	;
336	:	data_f1=	-494	;
337	:	data_f1=	493	;
338	:	data_f1=	1021	;
339	:	data_f1=	601	;
340	:	data_f1=	-377	;
341	:	data_f1=	-1006	;
342	:	data_f1=	-701	;
343	:	data_f1=	254	;
344	:	data_f1=	973	;
345	:	data_f1=	789	;
346	:	data_f1=	-129	;
347	:	data_f1=	-927	;
348	:	data_f1=	-865	;
349	:	data_f1=	0	;
350	:	data_f1=	864	;
351	:	data_f1=	926	;
352	:	data_f1=	128	;
353	:	data_f1=	-790	;
354	:	data_f1=	-974	;
355	:	data_f1=	-255	;
356	:	data_f1=	700	;
357	:	data_f1=	1005	;
358	:	data_f1=	376	;
359	:	data_f1=	-602	;
360	:	data_f1=	-1022	;
361	:	data_f1=	-494	;
362	:	data_f1=	493	;
363	:	data_f1=	1021	;
364	:	data_f1=	601	;
365	:	data_f1=	-377	;
366	:	data_f1=	-1006	;
367	:	data_f1=	-701	;
368	:	data_f1=	254	;
369	:	data_f1=	973	;
370	:	data_f1=	789	;
371	:	data_f1=	-129	;
372	:	data_f1=	-927	;
373	:	data_f1=	-865	;
374	:	data_f1=	0	;
375	:	data_f1=	864	;
376	:	data_f1=	926	;
377	:	data_f1=	128	;
378	:	data_f1=	-790	;
379	:	data_f1=	-974	;
380	:	data_f1=	-255	;
381	:	data_f1=	700	;
382	:	data_f1=	1005	;
383	:	data_f1=	376	;
384	:	data_f1=	-602	;
385	:	data_f1=	-1022	;
386	:	data_f1=	-494	;
387	:	data_f1=	493	;
388	:	data_f1=	1021	;
389	:	data_f1=	601	;
390	:	data_f1=	-377	;
391	:	data_f1=	-1006	;
392	:	data_f1=	-701	;
393	:	data_f1=	254	;
394	:	data_f1=	973	;
395	:	data_f1=	789	;
396	:	data_f1=	-129	;
397	:	data_f1=	-927	;
398	:	data_f1=	-865	;
399	:	data_f1=	-1	;
400	:	data_f1=	864	;
401	:	data_f1=	926	;
402	:	data_f1=	128	;
403	:	data_f1=	-790	;
404	:	data_f1=	-974	;
405	:	data_f1=	-255	;
406	:	data_f1=	700	;
407	:	data_f1=	1005	;
408	:	data_f1=	376	;
409	:	data_f1=	-602	;
410	:	data_f1=	-1022	;
411	:	data_f1=	-494	;
412	:	data_f1=	493	;
413	:	data_f1=	1021	;
414	:	data_f1=	601	;
415	:	data_f1=	-377	;
416	:	data_f1=	-1006	;
417	:	data_f1=	-701	;
418	:	data_f1=	254	;
419	:	data_f1=	973	;
420	:	data_f1=	789	;
421	:	data_f1=	-129	;
422	:	data_f1=	-927	;
423	:	data_f1=	-865	;
424	:	data_f1=	0	;
425	:	data_f1=	864	;
426	:	data_f1=	926	;
427	:	data_f1=	128	;
428	:	data_f1=	-790	;
429	:	data_f1=	-974	;
430	:	data_f1=	-255	;
431	:	data_f1=	700	;
432	:	data_f1=	1005	;
433	:	data_f1=	376	;
434	:	data_f1=	-602	;
435	:	data_f1=	-1022	;
436	:	data_f1=	-494	;
437	:	data_f1=	493	;
438	:	data_f1=	1021	;
439	:	data_f1=	601	;
440	:	data_f1=	-377	;
441	:	data_f1=	-1006	;
442	:	data_f1=	-701	;
443	:	data_f1=	254	;
444	:	data_f1=	973	;
445	:	data_f1=	789	;
446	:	data_f1=	-129	;
447	:	data_f1=	-927	;
448	:	data_f1=	-865	;
449	:	data_f1=	-1	;
450	:	data_f1=	864	;
451	:	data_f1=	926	;
452	:	data_f1=	128	;
453	:	data_f1=	-790	;
454	:	data_f1=	-974	;
455	:	data_f1=	-255	;
456	:	data_f1=	700	;
457	:	data_f1=	1005	;
458	:	data_f1=	376	;
459	:	data_f1=	-602	;
460	:	data_f1=	-1022	;
461	:	data_f1=	-494	;
462	:	data_f1=	493	;
463	:	data_f1=	1021	;
464	:	data_f1=	601	;
465	:	data_f1=	-377	;
466	:	data_f1=	-1006	;
467	:	data_f1=	-701	;
468	:	data_f1=	254	;
469	:	data_f1=	973	;
470	:	data_f1=	789	;
471	:	data_f1=	-129	;
472	:	data_f1=	-927	;
473	:	data_f1=	-865	;
474	:	data_f1=	-1	;
475	:	data_f1=	864	;
476	:	data_f1=	926	;
477	:	data_f1=	128	;
478	:	data_f1=	-790	;
479	:	data_f1=	-974	;
480	:	data_f1=	-255	;
481	:	data_f1=	700	;
482	:	data_f1=	1005	;
483	:	data_f1=	376	;
484	:	data_f1=	-602	;
485	:	data_f1=	-1022	;
486	:	data_f1=	-494	;
487	:	data_f1=	493	;
488	:	data_f1=	1021	;
489	:	data_f1=	601	;
490	:	data_f1=	-377	;
491	:	data_f1=	-1006	;
492	:	data_f1=	-701	;
493	:	data_f1=	254	;
494	:	data_f1=	973	;
495	:	data_f1=	789	;
496	:	data_f1=	-129	;
497	:	data_f1=	-927	;
498	:	data_f1=	-865	;
499	:	data_f1=	-1	;
500	:	data_f1=	864	;
501	:	data_f1=	926	;
502	:	data_f1=	128	;
503	:	data_f1=	-790	;
504	:	data_f1=	-974	;
505	:	data_f1=	-255	;
506	:	data_f1=	700	;
507	:	data_f1=	1005	;
508	:	data_f1=	376	;
509	:	data_f1=	-602	;
510	:	data_f1=	-1022	;
511	:	data_f1=	-494	;
512	:	data_f1=	493	;
513	:	data_f1=	1021	;
514	:	data_f1=	601	;
515	:	data_f1=	-377	;
516	:	data_f1=	-1006	;
517	:	data_f1=	-701	;
518	:	data_f1=	254	;
519	:	data_f1=	973	;
520	:	data_f1=	789	;
521	:	data_f1=	-129	;
522	:	data_f1=	-927	;
523	:	data_f1=	-865	;
524	:	data_f1=	0	;
525	:	data_f1=	864	;
526	:	data_f1=	926	;
527	:	data_f1=	128	;
528	:	data_f1=	-790	;
529	:	data_f1=	-974	;
530	:	data_f1=	-255	;
531	:	data_f1=	700	;
532	:	data_f1=	1005	;
533	:	data_f1=	376	;
534	:	data_f1=	-602	;
535	:	data_f1=	-1022	;
536	:	data_f1=	-494	;
537	:	data_f1=	493	;
538	:	data_f1=	1021	;
539	:	data_f1=	601	;
540	:	data_f1=	-377	;
541	:	data_f1=	-1006	;
542	:	data_f1=	-701	;
543	:	data_f1=	254	;
544	:	data_f1=	973	;
545	:	data_f1=	789	;
546	:	data_f1=	-129	;
547	:	data_f1=	-927	;
548	:	data_f1=	-865	;
549	:	data_f1=	-1	;
550	:	data_f1=	864	;
551	:	data_f1=	926	;
552	:	data_f1=	128	;
553	:	data_f1=	-790	;
554	:	data_f1=	-974	;
555	:	data_f1=	-255	;
556	:	data_f1=	700	;
557	:	data_f1=	1005	;
558	:	data_f1=	376	;
559	:	data_f1=	-602	;
560	:	data_f1=	-1022	;
561	:	data_f1=	-494	;
562	:	data_f1=	493	;
563	:	data_f1=	1021	;
564	:	data_f1=	601	;
565	:	data_f1=	-377	;
566	:	data_f1=	-1006	;
567	:	data_f1=	-701	;
568	:	data_f1=	254	;
569	:	data_f1=	973	;
570	:	data_f1=	789	;
571	:	data_f1=	-129	;
572	:	data_f1=	-927	;
573	:	data_f1=	-865	;
574	:	data_f1=	-1	;
575	:	data_f1=	864	;
576	:	data_f1=	926	;
577	:	data_f1=	128	;
578	:	data_f1=	-790	;
579	:	data_f1=	-974	;
580	:	data_f1=	-255	;
581	:	data_f1=	700	;
582	:	data_f1=	1005	;
583	:	data_f1=	376	;
584	:	data_f1=	-602	;
585	:	data_f1=	-1022	;
586	:	data_f1=	-494	;
587	:	data_f1=	493	;
588	:	data_f1=	1021	;
589	:	data_f1=	601	;
590	:	data_f1=	-377	;
591	:	data_f1=	-1006	;
592	:	data_f1=	-701	;
593	:	data_f1=	254	;
594	:	data_f1=	973	;
595	:	data_f1=	789	;
596	:	data_f1=	-129	;
597	:	data_f1=	-927	;
598	:	data_f1=	-865	;
599	:	data_f1=	-1	;
600	:	data_f1=	864	;
601	:	data_f1=	926	;
602	:	data_f1=	128	;
603	:	data_f1=	-790	;
604	:	data_f1=	-974	;
605	:	data_f1=	-255	;
606	:	data_f1=	700	;
607	:	data_f1=	1005	;
608	:	data_f1=	376	;
609	:	data_f1=	-602	;
610	:	data_f1=	-1022	;
611	:	data_f1=	-494	;
612	:	data_f1=	493	;
613	:	data_f1=	1021	;
614	:	data_f1=	601	;
615	:	data_f1=	-377	;
616	:	data_f1=	-1006	;
617	:	data_f1=	-701	;
618	:	data_f1=	254	;
619	:	data_f1=	973	;
620	:	data_f1=	789	;
621	:	data_f1=	-129	;
622	:	data_f1=	-927	;
623	:	data_f1=	-865	;
624	:	data_f1=	0	;
625	:	data_f1=	864	;
626	:	data_f1=	926	;
627	:	data_f1=	128	;
628	:	data_f1=	-790	;
629	:	data_f1=	-974	;
630	:	data_f1=	-255	;
631	:	data_f1=	700	;
632	:	data_f1=	1005	;
633	:	data_f1=	376	;
634	:	data_f1=	-602	;
635	:	data_f1=	-1022	;
636	:	data_f1=	-494	;
637	:	data_f1=	493	;
638	:	data_f1=	1021	;
639	:	data_f1=	601	;
640	:	data_f1=	-377	;
641	:	data_f1=	-1006	;
642	:	data_f1=	-701	;
643	:	data_f1=	254	;
644	:	data_f1=	973	;
645	:	data_f1=	789	;
646	:	data_f1=	-129	;
647	:	data_f1=	-927	;
648	:	data_f1=	-865	;
649	:	data_f1=	-1	;
650	:	data_f1=	864	;
651	:	data_f1=	926	;
652	:	data_f1=	128	;
653	:	data_f1=	-790	;
654	:	data_f1=	-974	;
655	:	data_f1=	-255	;
656	:	data_f1=	700	;
657	:	data_f1=	1005	;
658	:	data_f1=	376	;
659	:	data_f1=	-602	;
660	:	data_f1=	-1022	;
661	:	data_f1=	-494	;
662	:	data_f1=	493	;
663	:	data_f1=	1021	;
664	:	data_f1=	601	;
665	:	data_f1=	-377	;
666	:	data_f1=	-1006	;
667	:	data_f1=	-701	;
668	:	data_f1=	254	;
669	:	data_f1=	973	;
670	:	data_f1=	789	;
671	:	data_f1=	-129	;
672	:	data_f1=	-927	;
673	:	data_f1=	-865	;
674	:	data_f1=	-1	;
675	:	data_f1=	864	;
676	:	data_f1=	926	;
677	:	data_f1=	128	;
678	:	data_f1=	-790	;
679	:	data_f1=	-974	;
680	:	data_f1=	-255	;
681	:	data_f1=	700	;
682	:	data_f1=	1005	;
683	:	data_f1=	376	;
684	:	data_f1=	-602	;
685	:	data_f1=	-1022	;
686	:	data_f1=	-494	;
687	:	data_f1=	493	;
688	:	data_f1=	1021	;
689	:	data_f1=	601	;
690	:	data_f1=	-377	;
691	:	data_f1=	-1006	;
692	:	data_f1=	-701	;
693	:	data_f1=	254	;
694	:	data_f1=	973	;
695	:	data_f1=	789	;
696	:	data_f1=	-129	;
697	:	data_f1=	-927	;
698	:	data_f1=	-865	;
699	:	data_f1=	-1	;
700	:	data_f1=	864	;
701	:	data_f1=	926	;
702	:	data_f1=	128	;
703	:	data_f1=	-790	;
704	:	data_f1=	-974	;
705	:	data_f1=	-255	;
706	:	data_f1=	700	;
707	:	data_f1=	1005	;
708	:	data_f1=	376	;
709	:	data_f1=	-602	;
710	:	data_f1=	-1022	;
711	:	data_f1=	-494	;
712	:	data_f1=	493	;
713	:	data_f1=	1021	;
714	:	data_f1=	601	;
715	:	data_f1=	-377	;
716	:	data_f1=	-1006	;
717	:	data_f1=	-701	;
718	:	data_f1=	254	;
719	:	data_f1=	973	;
720	:	data_f1=	789	;
721	:	data_f1=	-129	;
722	:	data_f1=	-927	;
723	:	data_f1=	-865	;
724	:	data_f1=	0	;
725	:	data_f1=	864	;
726	:	data_f1=	926	;
727	:	data_f1=	128	;
728	:	data_f1=	-790	;
729	:	data_f1=	-974	;
730	:	data_f1=	-255	;
731	:	data_f1=	700	;
732	:	data_f1=	1005	;
733	:	data_f1=	376	;
734	:	data_f1=	-602	;
735	:	data_f1=	-1022	;
736	:	data_f1=	-494	;
737	:	data_f1=	493	;
738	:	data_f1=	1021	;
739	:	data_f1=	601	;
740	:	data_f1=	-377	;
741	:	data_f1=	-1006	;
742	:	data_f1=	-701	;
743	:	data_f1=	254	;
744	:	data_f1=	973	;
745	:	data_f1=	789	;
746	:	data_f1=	-129	;
747	:	data_f1=	-927	;
748	:	data_f1=	-865	;
749	:	data_f1=	0	;
750	:	data_f1=	864	;
751	:	data_f1=	926	;
752	:	data_f1=	128	;
753	:	data_f1=	-790	;
754	:	data_f1=	-974	;
755	:	data_f1=	-255	;
756	:	data_f1=	700	;
757	:	data_f1=	1005	;
758	:	data_f1=	376	;
759	:	data_f1=	-602	;
760	:	data_f1=	-1022	;
761	:	data_f1=	-494	;
762	:	data_f1=	493	;
763	:	data_f1=	1021	;
764	:	data_f1=	601	;
765	:	data_f1=	-377	;
766	:	data_f1=	-1006	;
767	:	data_f1=	-701	;
768	:	data_f1=	254	;
769	:	data_f1=	973	;
770	:	data_f1=	789	;
771	:	data_f1=	-129	;
772	:	data_f1=	-927	;
773	:	data_f1=	-865	;
774	:	data_f1=	-1	;
775	:	data_f1=	864	;
776	:	data_f1=	926	;
777	:	data_f1=	128	;
778	:	data_f1=	-790	;
779	:	data_f1=	-974	;
780	:	data_f1=	-255	;
781	:	data_f1=	700	;
782	:	data_f1=	1005	;
783	:	data_f1=	376	;
784	:	data_f1=	-602	;
785	:	data_f1=	-1022	;
786	:	data_f1=	-494	;
787	:	data_f1=	493	;
788	:	data_f1=	1021	;
789	:	data_f1=	601	;
790	:	data_f1=	-377	;
791	:	data_f1=	-1006	;
792	:	data_f1=	-701	;
793	:	data_f1=	254	;
794	:	data_f1=	973	;
795	:	data_f1=	789	;
796	:	data_f1=	-129	;
797	:	data_f1=	-927	;
798	:	data_f1=	-865	;
799	:	data_f1=	-1	;
800	:	data_f1=	864	;
801	:	data_f1=	926	;
802	:	data_f1=	128	;
803	:	data_f1=	-790	;
804	:	data_f1=	-974	;
805	:	data_f1=	-255	;
806	:	data_f1=	700	;
807	:	data_f1=	1005	;
808	:	data_f1=	376	;
809	:	data_f1=	-602	;
810	:	data_f1=	-1022	;
811	:	data_f1=	-494	;
812	:	data_f1=	493	;
813	:	data_f1=	1021	;
814	:	data_f1=	601	;
815	:	data_f1=	-377	;
816	:	data_f1=	-1006	;
817	:	data_f1=	-701	;
818	:	data_f1=	254	;
819	:	data_f1=	973	;
820	:	data_f1=	789	;
821	:	data_f1=	-129	;
822	:	data_f1=	-927	;
823	:	data_f1=	-865	;
824	:	data_f1=	-1	;
825	:	data_f1=	864	;
826	:	data_f1=	926	;
827	:	data_f1=	128	;
828	:	data_f1=	-790	;
829	:	data_f1=	-974	;
830	:	data_f1=	-255	;
831	:	data_f1=	700	;
832	:	data_f1=	1005	;
833	:	data_f1=	376	;
834	:	data_f1=	-602	;
835	:	data_f1=	-1022	;
836	:	data_f1=	-494	;
837	:	data_f1=	493	;
838	:	data_f1=	1021	;
839	:	data_f1=	601	;
840	:	data_f1=	-377	;
841	:	data_f1=	-1006	;
842	:	data_f1=	-701	;
843	:	data_f1=	254	;
844	:	data_f1=	973	;
845	:	data_f1=	789	;
846	:	data_f1=	-129	;
847	:	data_f1=	-927	;
848	:	data_f1=	-865	;
849	:	data_f1=	0	;
850	:	data_f1=	864	;
851	:	data_f1=	926	;
852	:	data_f1=	128	;
853	:	data_f1=	-790	;
854	:	data_f1=	-974	;
855	:	data_f1=	-255	;
856	:	data_f1=	700	;
857	:	data_f1=	1005	;
858	:	data_f1=	376	;
859	:	data_f1=	-602	;
860	:	data_f1=	-1022	;
861	:	data_f1=	-494	;
862	:	data_f1=	493	;
863	:	data_f1=	1021	;
864	:	data_f1=	601	;
865	:	data_f1=	-377	;
866	:	data_f1=	-1006	;
867	:	data_f1=	-701	;
868	:	data_f1=	254	;
869	:	data_f1=	973	;
870	:	data_f1=	789	;
871	:	data_f1=	-129	;
872	:	data_f1=	-927	;
873	:	data_f1=	-865	;
874	:	data_f1=	-1	;
875	:	data_f1=	864	;
876	:	data_f1=	926	;
877	:	data_f1=	128	;
878	:	data_f1=	-790	;
879	:	data_f1=	-974	;
880	:	data_f1=	-255	;
881	:	data_f1=	700	;
882	:	data_f1=	1005	;
883	:	data_f1=	376	;
884	:	data_f1=	-602	;
885	:	data_f1=	-1022	;
886	:	data_f1=	-494	;
887	:	data_f1=	493	;
888	:	data_f1=	1021	;
889	:	data_f1=	601	;
890	:	data_f1=	-377	;
891	:	data_f1=	-1006	;
892	:	data_f1=	-701	;
893	:	data_f1=	254	;
894	:	data_f1=	973	;
895	:	data_f1=	789	;
896	:	data_f1=	-129	;
897	:	data_f1=	-927	;
898	:	data_f1=	-865	;
899	:	data_f1=	-1	;
900	:	data_f1=	864	;
901	:	data_f1=	926	;
902	:	data_f1=	128	;
903	:	data_f1=	-790	;
904	:	data_f1=	-974	;
905	:	data_f1=	-255	;
906	:	data_f1=	700	;
907	:	data_f1=	1005	;
908	:	data_f1=	376	;
909	:	data_f1=	-602	;
910	:	data_f1=	-1022	;
911	:	data_f1=	-494	;
912	:	data_f1=	493	;
913	:	data_f1=	1021	;
914	:	data_f1=	601	;
915	:	data_f1=	-377	;
916	:	data_f1=	-1006	;
917	:	data_f1=	-701	;
918	:	data_f1=	254	;
919	:	data_f1=	973	;
920	:	data_f1=	789	;
921	:	data_f1=	-129	;
922	:	data_f1=	-927	;
923	:	data_f1=	-865	;
924	:	data_f1=	-1	;
925	:	data_f1=	864	;
926	:	data_f1=	926	;
927	:	data_f1=	128	;
928	:	data_f1=	-790	;
929	:	data_f1=	-974	;
930	:	data_f1=	-255	;
931	:	data_f1=	700	;
932	:	data_f1=	1005	;
933	:	data_f1=	376	;
934	:	data_f1=	-602	;
935	:	data_f1=	-1022	;
936	:	data_f1=	-494	;
937	:	data_f1=	493	;
938	:	data_f1=	1021	;
939	:	data_f1=	601	;
940	:	data_f1=	-377	;
941	:	data_f1=	-1006	;
942	:	data_f1=	-701	;
943	:	data_f1=	254	;
944	:	data_f1=	973	;
945	:	data_f1=	789	;
946	:	data_f1=	-129	;
947	:	data_f1=	-927	;
948	:	data_f1=	-865	;
949	:	data_f1=	-1	;
950	:	data_f1=	864	;
951	:	data_f1=	926	;
952	:	data_f1=	128	;
953	:	data_f1=	-790	;
954	:	data_f1=	-974	;
955	:	data_f1=	-255	;
956	:	data_f1=	700	;
957	:	data_f1=	1005	;
958	:	data_f1=	376	;
959	:	data_f1=	-602	;
960	:	data_f1=	-1022	;
961	:	data_f1=	-494	;
962	:	data_f1=	493	;
963	:	data_f1=	1021	;
964	:	data_f1=	601	;
965	:	data_f1=	-377	;
966	:	data_f1=	-1006	;
967	:	data_f1=	-701	;
968	:	data_f1=	254	;
969	:	data_f1=	973	;
970	:	data_f1=	789	;
971	:	data_f1=	-129	;
972	:	data_f1=	-927	;
973	:	data_f1=	-865	;
974	:	data_f1=	-1	;
975	:	data_f1=	864	;
976	:	data_f1=	926	;
977	:	data_f1=	128	;
978	:	data_f1=	-790	;
979	:	data_f1=	-974	;
980	:	data_f1=	-255	;
981	:	data_f1=	700	;
982	:	data_f1=	1005	;
983	:	data_f1=	376	;
984	:	data_f1=	-602	;
985	:	data_f1=	-1022	;
986	:	data_f1=	-494	;
987	:	data_f1=	493	;
988	:	data_f1=	1021	;
989	:	data_f1=	601	;
990	:	data_f1=	-377	;
991	:	data_f1=	-1006	;
992	:	data_f1=	-701	;
993	:	data_f1=	254	;
994	:	data_f1=	973	;
995	:	data_f1=	789	;
996	:	data_f1=	-129	;
997	:	data_f1=	-927	;
998	:	data_f1=	-865	;
999	:	data_f1=	-1	;
1000	:	data_f1=	0	;

default data_f1= 0;
endcase
always @*
case(count)
0	:	data_f2=	746	;
1	:	data_f2=	1021	;
2	:	data_f2=	652	;
3	:	data_f2=	-129	;
4	:	data_f2=	-829	;
5	:	data_f2=	-1006	;
6	:	data_f2=	-549	;
7	:	data_f2=	254	;
8	:	data_f2=	897	;
9	:	data_f2=	973	;
10	:	data_f2=	435	;
11	:	data_f2=	-377	;
12	:	data_f2=	-953	;
13	:	data_f2=	-927	;
14	:	data_f2=	-317	;
15	:	data_f2=	493	;
16	:	data_f2=	991	;
17	:	data_f2=	864	;
18	:	data_f2=	191	;
19	:	data_f2=	-602	;
20	:	data_f2=	-1016	;
21	:	data_f2=	-790	;
22	:	data_f2=	-65	;
23	:	data_f2=	700	;
24	:	data_f2=	1024	;
25	:	data_f2=	700	;
26	:	data_f2=	-65	;
27	:	data_f2=	-790	;
28	:	data_f2=	-1016	;
29	:	data_f2=	-602	;
30	:	data_f2=	191	;
31	:	data_f2=	864	;
32	:	data_f2=	991	;
33	:	data_f2=	493	;
34	:	data_f2=	-317	;
35	:	data_f2=	-927	;
36	:	data_f2=	-953	;
37	:	data_f2=	-377	;
38	:	data_f2=	435	;
39	:	data_f2=	973	;
40	:	data_f2=	897	;
41	:	data_f2=	254	;
42	:	data_f2=	-549	;
43	:	data_f2=	-1006	;
44	:	data_f2=	-829	;
45	:	data_f2=	-129	;
46	:	data_f2=	652	;
47	:	data_f2=	1021	;
48	:	data_f2=	746	;
49	:	data_f2=	-1	;
50	:	data_f2=	-747	;
51	:	data_f2=	-1022	;
52	:	data_f2=	-653	;
53	:	data_f2=	128	;
54	:	data_f2=	828	;
55	:	data_f2=	1005	;
56	:	data_f2=	548	;
57	:	data_f2=	-255	;
58	:	data_f2=	-898	;
59	:	data_f2=	-974	;
60	:	data_f2=	-436	;
61	:	data_f2=	376	;
62	:	data_f2=	952	;
63	:	data_f2=	926	;
64	:	data_f2=	316	;
65	:	data_f2=	-494	;
66	:	data_f2=	-992	;
67	:	data_f2=	-865	;
68	:	data_f2=	-192	;
69	:	data_f2=	601	;
70	:	data_f2=	1015	;
71	:	data_f2=	789	;
72	:	data_f2=	64	;
73	:	data_f2=	-701	;
74	:	data_f2=	-1024	;
75	:	data_f2=	-701	;
76	:	data_f2=	64	;
77	:	data_f2=	789	;
78	:	data_f2=	1015	;
79	:	data_f2=	601	;
80	:	data_f2=	-192	;
81	:	data_f2=	-865	;
82	:	data_f2=	-992	;
83	:	data_f2=	-494	;
84	:	data_f2=	316	;
85	:	data_f2=	926	;
86	:	data_f2=	952	;
87	:	data_f2=	376	;
88	:	data_f2=	-436	;
89	:	data_f2=	-974	;
90	:	data_f2=	-898	;
91	:	data_f2=	-255	;
92	:	data_f2=	548	;
93	:	data_f2=	1005	;
94	:	data_f2=	828	;
95	:	data_f2=	128	;
96	:	data_f2=	-653	;
97	:	data_f2=	-1022	;
98	:	data_f2=	-747	;
99	:	data_f2=	0	;
100	:	data_f2=	746	;
101	:	data_f2=	1021	;
102	:	data_f2=	652	;
103	:	data_f2=	-129	;
104	:	data_f2=	-829	;
105	:	data_f2=	-1006	;
106	:	data_f2=	-549	;
107	:	data_f2=	254	;
108	:	data_f2=	897	;
109	:	data_f2=	973	;
110	:	data_f2=	435	;
111	:	data_f2=	-377	;
112	:	data_f2=	-953	;
113	:	data_f2=	-927	;
114	:	data_f2=	-317	;
115	:	data_f2=	493	;
116	:	data_f2=	991	;
117	:	data_f2=	864	;
118	:	data_f2=	191	;
119	:	data_f2=	-602	;
120	:	data_f2=	-1016	;
121	:	data_f2=	-790	;
122	:	data_f2=	-65	;
123	:	data_f2=	700	;
124	:	data_f2=	1024	;
125	:	data_f2=	700	;
126	:	data_f2=	-65	;
127	:	data_f2=	-790	;
128	:	data_f2=	-1016	;
129	:	data_f2=	-602	;
130	:	data_f2=	191	;
131	:	data_f2=	864	;
132	:	data_f2=	991	;
133	:	data_f2=	493	;
134	:	data_f2=	-317	;
135	:	data_f2=	-927	;
136	:	data_f2=	-953	;
137	:	data_f2=	-377	;
138	:	data_f2=	435	;
139	:	data_f2=	973	;
140	:	data_f2=	897	;
141	:	data_f2=	254	;
142	:	data_f2=	-549	;
143	:	data_f2=	-1006	;
144	:	data_f2=	-829	;
145	:	data_f2=	-129	;
146	:	data_f2=	652	;
147	:	data_f2=	1021	;
148	:	data_f2=	746	;
149	:	data_f2=	-1	;
150	:	data_f2=	-747	;
151	:	data_f2=	-1022	;
152	:	data_f2=	-653	;
153	:	data_f2=	128	;
154	:	data_f2=	828	;
155	:	data_f2=	1005	;
156	:	data_f2=	548	;
157	:	data_f2=	-255	;
158	:	data_f2=	-898	;
159	:	data_f2=	-974	;
160	:	data_f2=	-436	;
161	:	data_f2=	376	;
162	:	data_f2=	952	;
163	:	data_f2=	926	;
164	:	data_f2=	316	;
165	:	data_f2=	-494	;
166	:	data_f2=	-992	;
167	:	data_f2=	-865	;
168	:	data_f2=	-192	;
169	:	data_f2=	601	;
170	:	data_f2=	1015	;
171	:	data_f2=	789	;
172	:	data_f2=	64	;
173	:	data_f2=	-701	;
174	:	data_f2=	-1024	;
175	:	data_f2=	-701	;
176	:	data_f2=	64	;
177	:	data_f2=	789	;
178	:	data_f2=	1015	;
179	:	data_f2=	601	;
180	:	data_f2=	-192	;
181	:	data_f2=	-865	;
182	:	data_f2=	-992	;
183	:	data_f2=	-494	;
184	:	data_f2=	316	;
185	:	data_f2=	926	;
186	:	data_f2=	952	;
187	:	data_f2=	376	;
188	:	data_f2=	-436	;
189	:	data_f2=	-974	;
190	:	data_f2=	-898	;
191	:	data_f2=	-255	;
192	:	data_f2=	548	;
193	:	data_f2=	1005	;
194	:	data_f2=	828	;
195	:	data_f2=	128	;
196	:	data_f2=	-653	;
197	:	data_f2=	-1022	;
198	:	data_f2=	-747	;
199	:	data_f2=	0	;
200	:	data_f2=	746	;
201	:	data_f2=	1021	;
202	:	data_f2=	652	;
203	:	data_f2=	-129	;
204	:	data_f2=	-829	;
205	:	data_f2=	-1006	;
206	:	data_f2=	-549	;
207	:	data_f2=	254	;
208	:	data_f2=	897	;
209	:	data_f2=	973	;
210	:	data_f2=	435	;
211	:	data_f2=	-377	;
212	:	data_f2=	-953	;
213	:	data_f2=	-927	;
214	:	data_f2=	-317	;
215	:	data_f2=	493	;
216	:	data_f2=	991	;
217	:	data_f2=	864	;
218	:	data_f2=	191	;
219	:	data_f2=	-602	;
220	:	data_f2=	-1016	;
221	:	data_f2=	-790	;
222	:	data_f2=	-65	;
223	:	data_f2=	700	;
224	:	data_f2=	1024	;
225	:	data_f2=	700	;
226	:	data_f2=	-65	;
227	:	data_f2=	-790	;
228	:	data_f2=	-1016	;
229	:	data_f2=	-602	;
230	:	data_f2=	191	;
231	:	data_f2=	864	;
232	:	data_f2=	991	;
233	:	data_f2=	493	;
234	:	data_f2=	-317	;
235	:	data_f2=	-927	;
236	:	data_f2=	-953	;
237	:	data_f2=	-377	;
238	:	data_f2=	435	;
239	:	data_f2=	973	;
240	:	data_f2=	897	;
241	:	data_f2=	254	;
242	:	data_f2=	-549	;
243	:	data_f2=	-1006	;
244	:	data_f2=	-829	;
245	:	data_f2=	-129	;
246	:	data_f2=	652	;
247	:	data_f2=	1021	;
248	:	data_f2=	746	;
249	:	data_f2=	-1	;
250	:	data_f2=	-747	;
251	:	data_f2=	-1022	;
252	:	data_f2=	-653	;
253	:	data_f2=	128	;
254	:	data_f2=	828	;
255	:	data_f2=	1005	;
256	:	data_f2=	548	;
257	:	data_f2=	-255	;
258	:	data_f2=	-898	;
259	:	data_f2=	-974	;
260	:	data_f2=	-436	;
261	:	data_f2=	376	;
262	:	data_f2=	952	;
263	:	data_f2=	926	;
264	:	data_f2=	316	;
265	:	data_f2=	-494	;
266	:	data_f2=	-992	;
267	:	data_f2=	-865	;
268	:	data_f2=	-192	;
269	:	data_f2=	601	;
270	:	data_f2=	1015	;
271	:	data_f2=	789	;
272	:	data_f2=	64	;
273	:	data_f2=	-701	;
274	:	data_f2=	-1024	;
275	:	data_f2=	-701	;
276	:	data_f2=	64	;
277	:	data_f2=	789	;
278	:	data_f2=	1015	;
279	:	data_f2=	601	;
280	:	data_f2=	-192	;
281	:	data_f2=	-865	;
282	:	data_f2=	-992	;
283	:	data_f2=	-494	;
284	:	data_f2=	316	;
285	:	data_f2=	926	;
286	:	data_f2=	952	;
287	:	data_f2=	376	;
288	:	data_f2=	-436	;
289	:	data_f2=	-974	;
290	:	data_f2=	-898	;
291	:	data_f2=	-255	;
292	:	data_f2=	548	;
293	:	data_f2=	1005	;
294	:	data_f2=	828	;
295	:	data_f2=	128	;
296	:	data_f2=	-653	;
297	:	data_f2=	-1022	;
298	:	data_f2=	-747	;
299	:	data_f2=	0	;
300	:	data_f2=	746	;
301	:	data_f2=	1021	;
302	:	data_f2=	652	;
303	:	data_f2=	-129	;
304	:	data_f2=	-829	;
305	:	data_f2=	-1006	;
306	:	data_f2=	-549	;
307	:	data_f2=	254	;
308	:	data_f2=	897	;
309	:	data_f2=	973	;
310	:	data_f2=	435	;
311	:	data_f2=	-377	;
312	:	data_f2=	-953	;
313	:	data_f2=	-927	;
314	:	data_f2=	-317	;
315	:	data_f2=	493	;
316	:	data_f2=	991	;
317	:	data_f2=	864	;
318	:	data_f2=	191	;
319	:	data_f2=	-602	;
320	:	data_f2=	-1016	;
321	:	data_f2=	-790	;
322	:	data_f2=	-65	;
323	:	data_f2=	700	;
324	:	data_f2=	1024	;
325	:	data_f2=	700	;
326	:	data_f2=	-65	;
327	:	data_f2=	-790	;
328	:	data_f2=	-1016	;
329	:	data_f2=	-602	;
330	:	data_f2=	191	;
331	:	data_f2=	864	;
332	:	data_f2=	991	;
333	:	data_f2=	493	;
334	:	data_f2=	-317	;
335	:	data_f2=	-927	;
336	:	data_f2=	-953	;
337	:	data_f2=	-377	;
338	:	data_f2=	435	;
339	:	data_f2=	973	;
340	:	data_f2=	897	;
341	:	data_f2=	254	;
342	:	data_f2=	-549	;
343	:	data_f2=	-1006	;
344	:	data_f2=	-829	;
345	:	data_f2=	-129	;
346	:	data_f2=	652	;
347	:	data_f2=	1021	;
348	:	data_f2=	746	;
349	:	data_f2=	-1	;
350	:	data_f2=	-747	;
351	:	data_f2=	-1022	;
352	:	data_f2=	-653	;
353	:	data_f2=	128	;
354	:	data_f2=	828	;
355	:	data_f2=	1005	;
356	:	data_f2=	548	;
357	:	data_f2=	-255	;
358	:	data_f2=	-898	;
359	:	data_f2=	-974	;
360	:	data_f2=	-436	;
361	:	data_f2=	376	;
362	:	data_f2=	952	;
363	:	data_f2=	926	;
364	:	data_f2=	316	;
365	:	data_f2=	-494	;
366	:	data_f2=	-992	;
367	:	data_f2=	-865	;
368	:	data_f2=	-192	;
369	:	data_f2=	601	;
370	:	data_f2=	1015	;
371	:	data_f2=	789	;
372	:	data_f2=	64	;
373	:	data_f2=	-701	;
374	:	data_f2=	-1024	;
375	:	data_f2=	-701	;
376	:	data_f2=	64	;
377	:	data_f2=	789	;
378	:	data_f2=	1015	;
379	:	data_f2=	601	;
380	:	data_f2=	-192	;
381	:	data_f2=	-865	;
382	:	data_f2=	-992	;
383	:	data_f2=	-494	;
384	:	data_f2=	316	;
385	:	data_f2=	926	;
386	:	data_f2=	952	;
387	:	data_f2=	376	;
388	:	data_f2=	-436	;
389	:	data_f2=	-974	;
390	:	data_f2=	-898	;
391	:	data_f2=	-255	;
392	:	data_f2=	548	;
393	:	data_f2=	1005	;
394	:	data_f2=	828	;
395	:	data_f2=	128	;
396	:	data_f2=	-653	;
397	:	data_f2=	-1022	;
398	:	data_f2=	-747	;
399	:	data_f2=	0	;
400	:	data_f2=	746	;
401	:	data_f2=	1021	;
402	:	data_f2=	652	;
403	:	data_f2=	-129	;
404	:	data_f2=	-829	;
405	:	data_f2=	-1006	;
406	:	data_f2=	-549	;
407	:	data_f2=	254	;
408	:	data_f2=	897	;
409	:	data_f2=	973	;
410	:	data_f2=	435	;
411	:	data_f2=	-377	;
412	:	data_f2=	-953	;
413	:	data_f2=	-927	;
414	:	data_f2=	-317	;
415	:	data_f2=	493	;
416	:	data_f2=	991	;
417	:	data_f2=	864	;
418	:	data_f2=	191	;
419	:	data_f2=	-602	;
420	:	data_f2=	-1016	;
421	:	data_f2=	-790	;
422	:	data_f2=	-65	;
423	:	data_f2=	700	;
424	:	data_f2=	1024	;
425	:	data_f2=	700	;
426	:	data_f2=	-65	;
427	:	data_f2=	-790	;
428	:	data_f2=	-1016	;
429	:	data_f2=	-602	;
430	:	data_f2=	191	;
431	:	data_f2=	864	;
432	:	data_f2=	991	;
433	:	data_f2=	493	;
434	:	data_f2=	-317	;
435	:	data_f2=	-927	;
436	:	data_f2=	-953	;
437	:	data_f2=	-377	;
438	:	data_f2=	435	;
439	:	data_f2=	973	;
440	:	data_f2=	897	;
441	:	data_f2=	254	;
442	:	data_f2=	-549	;
443	:	data_f2=	-1006	;
444	:	data_f2=	-829	;
445	:	data_f2=	-129	;
446	:	data_f2=	652	;
447	:	data_f2=	1021	;
448	:	data_f2=	746	;
449	:	data_f2=	0	;
450	:	data_f2=	-747	;
451	:	data_f2=	-1022	;
452	:	data_f2=	-653	;
453	:	data_f2=	128	;
454	:	data_f2=	828	;
455	:	data_f2=	1005	;
456	:	data_f2=	548	;
457	:	data_f2=	-255	;
458	:	data_f2=	-898	;
459	:	data_f2=	-974	;
460	:	data_f2=	-436	;
461	:	data_f2=	376	;
462	:	data_f2=	952	;
463	:	data_f2=	926	;
464	:	data_f2=	316	;
465	:	data_f2=	-494	;
466	:	data_f2=	-992	;
467	:	data_f2=	-865	;
468	:	data_f2=	-192	;
469	:	data_f2=	601	;
470	:	data_f2=	1015	;
471	:	data_f2=	789	;
472	:	data_f2=	64	;
473	:	data_f2=	-701	;
474	:	data_f2=	-1024	;
475	:	data_f2=	-701	;
476	:	data_f2=	64	;
477	:	data_f2=	789	;
478	:	data_f2=	1015	;
479	:	data_f2=	601	;
480	:	data_f2=	-192	;
481	:	data_f2=	-865	;
482	:	data_f2=	-992	;
483	:	data_f2=	-494	;
484	:	data_f2=	316	;
485	:	data_f2=	926	;
486	:	data_f2=	952	;
487	:	data_f2=	376	;
488	:	data_f2=	-436	;
489	:	data_f2=	-974	;
490	:	data_f2=	-898	;
491	:	data_f2=	-255	;
492	:	data_f2=	548	;
493	:	data_f2=	1005	;
494	:	data_f2=	828	;
495	:	data_f2=	128	;
496	:	data_f2=	-653	;
497	:	data_f2=	-1022	;
498	:	data_f2=	-747	;
499	:	data_f2=	0	;
500	:	data_f2=	746	;
501	:	data_f2=	1021	;
502	:	data_f2=	652	;
503	:	data_f2=	-129	;
504	:	data_f2=	-829	;
505	:	data_f2=	-1006	;
506	:	data_f2=	-549	;
507	:	data_f2=	254	;
508	:	data_f2=	897	;
509	:	data_f2=	973	;
510	:	data_f2=	435	;
511	:	data_f2=	-377	;
512	:	data_f2=	-953	;
513	:	data_f2=	-927	;
514	:	data_f2=	-317	;
515	:	data_f2=	493	;
516	:	data_f2=	991	;
517	:	data_f2=	864	;
518	:	data_f2=	191	;
519	:	data_f2=	-602	;
520	:	data_f2=	-1016	;
521	:	data_f2=	-790	;
522	:	data_f2=	-65	;
523	:	data_f2=	700	;
524	:	data_f2=	1024	;
525	:	data_f2=	700	;
526	:	data_f2=	-65	;
527	:	data_f2=	-790	;
528	:	data_f2=	-1016	;
529	:	data_f2=	-602	;
530	:	data_f2=	191	;
531	:	data_f2=	864	;
532	:	data_f2=	991	;
533	:	data_f2=	493	;
534	:	data_f2=	-317	;
535	:	data_f2=	-927	;
536	:	data_f2=	-953	;
537	:	data_f2=	-377	;
538	:	data_f2=	435	;
539	:	data_f2=	973	;
540	:	data_f2=	897	;
541	:	data_f2=	254	;
542	:	data_f2=	-549	;
543	:	data_f2=	-1006	;
544	:	data_f2=	-829	;
545	:	data_f2=	-129	;
546	:	data_f2=	652	;
547	:	data_f2=	1021	;
548	:	data_f2=	746	;
549	:	data_f2=	0	;
550	:	data_f2=	-747	;
551	:	data_f2=	-1022	;
552	:	data_f2=	-653	;
553	:	data_f2=	128	;
554	:	data_f2=	828	;
555	:	data_f2=	1005	;
556	:	data_f2=	548	;
557	:	data_f2=	-255	;
558	:	data_f2=	-898	;
559	:	data_f2=	-974	;
560	:	data_f2=	-436	;
561	:	data_f2=	376	;
562	:	data_f2=	952	;
563	:	data_f2=	926	;
564	:	data_f2=	316	;
565	:	data_f2=	-494	;
566	:	data_f2=	-992	;
567	:	data_f2=	-865	;
568	:	data_f2=	-192	;
569	:	data_f2=	601	;
570	:	data_f2=	1015	;
571	:	data_f2=	789	;
572	:	data_f2=	64	;
573	:	data_f2=	-701	;
574	:	data_f2=	-1024	;
575	:	data_f2=	-701	;
576	:	data_f2=	64	;
577	:	data_f2=	789	;
578	:	data_f2=	1015	;
579	:	data_f2=	601	;
580	:	data_f2=	-192	;
581	:	data_f2=	-865	;
582	:	data_f2=	-992	;
583	:	data_f2=	-494	;
584	:	data_f2=	316	;
585	:	data_f2=	926	;
586	:	data_f2=	952	;
587	:	data_f2=	376	;
588	:	data_f2=	-436	;
589	:	data_f2=	-974	;
590	:	data_f2=	-898	;
591	:	data_f2=	-255	;
592	:	data_f2=	548	;
593	:	data_f2=	1005	;
594	:	data_f2=	828	;
595	:	data_f2=	128	;
596	:	data_f2=	-653	;
597	:	data_f2=	-1022	;
598	:	data_f2=	-747	;
599	:	data_f2=	0	;
600	:	data_f2=	746	;
601	:	data_f2=	1021	;
602	:	data_f2=	652	;
603	:	data_f2=	-129	;
604	:	data_f2=	-829	;
605	:	data_f2=	-1006	;
606	:	data_f2=	-549	;
607	:	data_f2=	254	;
608	:	data_f2=	897	;
609	:	data_f2=	973	;
610	:	data_f2=	435	;
611	:	data_f2=	-377	;
612	:	data_f2=	-953	;
613	:	data_f2=	-927	;
614	:	data_f2=	-317	;
615	:	data_f2=	493	;
616	:	data_f2=	991	;
617	:	data_f2=	864	;
618	:	data_f2=	191	;
619	:	data_f2=	-602	;
620	:	data_f2=	-1016	;
621	:	data_f2=	-790	;
622	:	data_f2=	-65	;
623	:	data_f2=	700	;
624	:	data_f2=	1024	;
625	:	data_f2=	700	;
626	:	data_f2=	-65	;
627	:	data_f2=	-790	;
628	:	data_f2=	-1016	;
629	:	data_f2=	-602	;
630	:	data_f2=	191	;
631	:	data_f2=	864	;
632	:	data_f2=	991	;
633	:	data_f2=	493	;
634	:	data_f2=	-317	;
635	:	data_f2=	-927	;
636	:	data_f2=	-953	;
637	:	data_f2=	-377	;
638	:	data_f2=	435	;
639	:	data_f2=	973	;
640	:	data_f2=	897	;
641	:	data_f2=	254	;
642	:	data_f2=	-549	;
643	:	data_f2=	-1006	;
644	:	data_f2=	-829	;
645	:	data_f2=	-129	;
646	:	data_f2=	652	;
647	:	data_f2=	1021	;
648	:	data_f2=	746	;
649	:	data_f2=	0	;
650	:	data_f2=	-747	;
651	:	data_f2=	-1022	;
652	:	data_f2=	-653	;
653	:	data_f2=	128	;
654	:	data_f2=	828	;
655	:	data_f2=	1005	;
656	:	data_f2=	548	;
657	:	data_f2=	-255	;
658	:	data_f2=	-898	;
659	:	data_f2=	-974	;
660	:	data_f2=	-436	;
661	:	data_f2=	376	;
662	:	data_f2=	952	;
663	:	data_f2=	926	;
664	:	data_f2=	316	;
665	:	data_f2=	-494	;
666	:	data_f2=	-992	;
667	:	data_f2=	-865	;
668	:	data_f2=	-192	;
669	:	data_f2=	601	;
670	:	data_f2=	1015	;
671	:	data_f2=	789	;
672	:	data_f2=	64	;
673	:	data_f2=	-701	;
674	:	data_f2=	-1024	;
675	:	data_f2=	-701	;
676	:	data_f2=	64	;
677	:	data_f2=	789	;
678	:	data_f2=	1015	;
679	:	data_f2=	601	;
680	:	data_f2=	-192	;
681	:	data_f2=	-865	;
682	:	data_f2=	-992	;
683	:	data_f2=	-494	;
684	:	data_f2=	316	;
685	:	data_f2=	926	;
686	:	data_f2=	952	;
687	:	data_f2=	376	;
688	:	data_f2=	-436	;
689	:	data_f2=	-974	;
690	:	data_f2=	-898	;
691	:	data_f2=	-255	;
692	:	data_f2=	548	;
693	:	data_f2=	1005	;
694	:	data_f2=	828	;
695	:	data_f2=	128	;
696	:	data_f2=	-653	;
697	:	data_f2=	-1022	;
698	:	data_f2=	-747	;
699	:	data_f2=	-1	;
700	:	data_f2=	746	;
701	:	data_f2=	1021	;
702	:	data_f2=	652	;
703	:	data_f2=	-129	;
704	:	data_f2=	-829	;
705	:	data_f2=	-1006	;
706	:	data_f2=	-549	;
707	:	data_f2=	254	;
708	:	data_f2=	897	;
709	:	data_f2=	973	;
710	:	data_f2=	435	;
711	:	data_f2=	-377	;
712	:	data_f2=	-953	;
713	:	data_f2=	-927	;
714	:	data_f2=	-317	;
715	:	data_f2=	493	;
716	:	data_f2=	991	;
717	:	data_f2=	864	;
718	:	data_f2=	191	;
719	:	data_f2=	-602	;
720	:	data_f2=	-1016	;
721	:	data_f2=	-790	;
722	:	data_f2=	-65	;
723	:	data_f2=	700	;
724	:	data_f2=	1024	;
725	:	data_f2=	700	;
726	:	data_f2=	-65	;
727	:	data_f2=	-790	;
728	:	data_f2=	-1016	;
729	:	data_f2=	-602	;
730	:	data_f2=	191	;
731	:	data_f2=	864	;
732	:	data_f2=	991	;
733	:	data_f2=	493	;
734	:	data_f2=	-317	;
735	:	data_f2=	-927	;
736	:	data_f2=	-953	;
737	:	data_f2=	-377	;
738	:	data_f2=	435	;
739	:	data_f2=	973	;
740	:	data_f2=	897	;
741	:	data_f2=	254	;
742	:	data_f2=	-549	;
743	:	data_f2=	-1006	;
744	:	data_f2=	-829	;
745	:	data_f2=	-129	;
746	:	data_f2=	652	;
747	:	data_f2=	1021	;
748	:	data_f2=	746	;
749	:	data_f2=	-1	;
750	:	data_f2=	-747	;
751	:	data_f2=	-1022	;
752	:	data_f2=	-653	;
753	:	data_f2=	128	;
754	:	data_f2=	828	;
755	:	data_f2=	1005	;
756	:	data_f2=	548	;
757	:	data_f2=	-255	;
758	:	data_f2=	-898	;
759	:	data_f2=	-974	;
760	:	data_f2=	-436	;
761	:	data_f2=	376	;
762	:	data_f2=	952	;
763	:	data_f2=	926	;
764	:	data_f2=	316	;
765	:	data_f2=	-494	;
766	:	data_f2=	-992	;
767	:	data_f2=	-865	;
768	:	data_f2=	-192	;
769	:	data_f2=	601	;
770	:	data_f2=	1015	;
771	:	data_f2=	789	;
772	:	data_f2=	64	;
773	:	data_f2=	-701	;
774	:	data_f2=	-1024	;
775	:	data_f2=	-701	;
776	:	data_f2=	64	;
777	:	data_f2=	789	;
778	:	data_f2=	1015	;
779	:	data_f2=	601	;
780	:	data_f2=	-192	;
781	:	data_f2=	-865	;
782	:	data_f2=	-992	;
783	:	data_f2=	-494	;
784	:	data_f2=	316	;
785	:	data_f2=	926	;
786	:	data_f2=	952	;
787	:	data_f2=	376	;
788	:	data_f2=	-436	;
789	:	data_f2=	-974	;
790	:	data_f2=	-898	;
791	:	data_f2=	-255	;
792	:	data_f2=	548	;
793	:	data_f2=	1005	;
794	:	data_f2=	828	;
795	:	data_f2=	128	;
796	:	data_f2=	-653	;
797	:	data_f2=	-1022	;
798	:	data_f2=	-747	;
799	:	data_f2=	0	;
800	:	data_f2=	746	;
801	:	data_f2=	1021	;
802	:	data_f2=	652	;
803	:	data_f2=	-129	;
804	:	data_f2=	-829	;
805	:	data_f2=	-1006	;
806	:	data_f2=	-549	;
807	:	data_f2=	254	;
808	:	data_f2=	897	;
809	:	data_f2=	973	;
810	:	data_f2=	435	;
811	:	data_f2=	-377	;
812	:	data_f2=	-953	;
813	:	data_f2=	-927	;
814	:	data_f2=	-317	;
815	:	data_f2=	493	;
816	:	data_f2=	991	;
817	:	data_f2=	864	;
818	:	data_f2=	191	;
819	:	data_f2=	-602	;
820	:	data_f2=	-1016	;
821	:	data_f2=	-790	;
822	:	data_f2=	-65	;
823	:	data_f2=	700	;
824	:	data_f2=	1024	;
825	:	data_f2=	700	;
826	:	data_f2=	-65	;
827	:	data_f2=	-790	;
828	:	data_f2=	-1016	;
829	:	data_f2=	-602	;
830	:	data_f2=	191	;
831	:	data_f2=	864	;
832	:	data_f2=	991	;
833	:	data_f2=	493	;
834	:	data_f2=	-317	;
835	:	data_f2=	-927	;
836	:	data_f2=	-953	;
837	:	data_f2=	-377	;
838	:	data_f2=	435	;
839	:	data_f2=	973	;
840	:	data_f2=	897	;
841	:	data_f2=	254	;
842	:	data_f2=	-549	;
843	:	data_f2=	-1006	;
844	:	data_f2=	-829	;
845	:	data_f2=	-129	;
846	:	data_f2=	652	;
847	:	data_f2=	1021	;
848	:	data_f2=	746	;
849	:	data_f2=	-1	;
850	:	data_f2=	-747	;
851	:	data_f2=	-1022	;
852	:	data_f2=	-653	;
853	:	data_f2=	128	;
854	:	data_f2=	828	;
855	:	data_f2=	1005	;
856	:	data_f2=	548	;
857	:	data_f2=	-255	;
858	:	data_f2=	-898	;
859	:	data_f2=	-974	;
860	:	data_f2=	-436	;
861	:	data_f2=	376	;
862	:	data_f2=	952	;
863	:	data_f2=	926	;
864	:	data_f2=	316	;
865	:	data_f2=	-494	;
866	:	data_f2=	-992	;
867	:	data_f2=	-865	;
868	:	data_f2=	-192	;
869	:	data_f2=	601	;
870	:	data_f2=	1015	;
871	:	data_f2=	789	;
872	:	data_f2=	64	;
873	:	data_f2=	-701	;
874	:	data_f2=	-1024	;
875	:	data_f2=	-701	;
876	:	data_f2=	64	;
877	:	data_f2=	789	;
878	:	data_f2=	1015	;
879	:	data_f2=	601	;
880	:	data_f2=	-192	;
881	:	data_f2=	-865	;
882	:	data_f2=	-992	;
883	:	data_f2=	-494	;
884	:	data_f2=	316	;
885	:	data_f2=	926	;
886	:	data_f2=	952	;
887	:	data_f2=	376	;
888	:	data_f2=	-436	;
889	:	data_f2=	-974	;
890	:	data_f2=	-898	;
891	:	data_f2=	-255	;
892	:	data_f2=	548	;
893	:	data_f2=	1005	;
894	:	data_f2=	828	;
895	:	data_f2=	128	;
896	:	data_f2=	-653	;
897	:	data_f2=	-1022	;
898	:	data_f2=	-747	;
899	:	data_f2=	0	;
900	:	data_f2=	746	;
901	:	data_f2=	1021	;
902	:	data_f2=	652	;
903	:	data_f2=	-129	;
904	:	data_f2=	-829	;
905	:	data_f2=	-1006	;
906	:	data_f2=	-549	;
907	:	data_f2=	254	;
908	:	data_f2=	897	;
909	:	data_f2=	973	;
910	:	data_f2=	435	;
911	:	data_f2=	-377	;
912	:	data_f2=	-953	;
913	:	data_f2=	-927	;
914	:	data_f2=	-317	;
915	:	data_f2=	493	;
916	:	data_f2=	991	;
917	:	data_f2=	864	;
918	:	data_f2=	191	;
919	:	data_f2=	-602	;
920	:	data_f2=	-1016	;
921	:	data_f2=	-790	;
922	:	data_f2=	-65	;
923	:	data_f2=	700	;
924	:	data_f2=	1024	;
925	:	data_f2=	700	;
926	:	data_f2=	-65	;
927	:	data_f2=	-790	;
928	:	data_f2=	-1016	;
929	:	data_f2=	-602	;
930	:	data_f2=	191	;
931	:	data_f2=	864	;
932	:	data_f2=	991	;
933	:	data_f2=	493	;
934	:	data_f2=	-317	;
935	:	data_f2=	-927	;
936	:	data_f2=	-953	;
937	:	data_f2=	-377	;
938	:	data_f2=	435	;
939	:	data_f2=	973	;
940	:	data_f2=	897	;
941	:	data_f2=	254	;
942	:	data_f2=	-549	;
943	:	data_f2=	-1006	;
944	:	data_f2=	-829	;
945	:	data_f2=	-129	;
946	:	data_f2=	652	;
947	:	data_f2=	1021	;
948	:	data_f2=	746	;
949	:	data_f2=	0	;
950	:	data_f2=	-747	;
951	:	data_f2=	-1022	;
952	:	data_f2=	-653	;
953	:	data_f2=	128	;
954	:	data_f2=	828	;
955	:	data_f2=	1005	;
956	:	data_f2=	548	;
957	:	data_f2=	-255	;
958	:	data_f2=	-898	;
959	:	data_f2=	-974	;
960	:	data_f2=	-436	;
961	:	data_f2=	376	;
962	:	data_f2=	952	;
963	:	data_f2=	926	;
964	:	data_f2=	316	;
965	:	data_f2=	-494	;
966	:	data_f2=	-992	;
967	:	data_f2=	-865	;
968	:	data_f2=	-192	;
969	:	data_f2=	601	;
970	:	data_f2=	1015	;
971	:	data_f2=	789	;
972	:	data_f2=	64	;
973	:	data_f2=	-701	;
974	:	data_f2=	-1024	;
975	:	data_f2=	-701	;
976	:	data_f2=	64	;
977	:	data_f2=	789	;
978	:	data_f2=	1015	;
979	:	data_f2=	601	;
980	:	data_f2=	-192	;
981	:	data_f2=	-865	;
982	:	data_f2=	-992	;
983	:	data_f2=	-494	;
984	:	data_f2=	316	;
985	:	data_f2=	926	;
986	:	data_f2=	952	;
987	:	data_f2=	376	;
988	:	data_f2=	-436	;
989	:	data_f2=	-974	;
990	:	data_f2=	-898	;
991	:	data_f2=	-255	;
992	:	data_f2=	548	;
993	:	data_f2=	1005	;
994	:	data_f2=	828	;
995	:	data_f2=	128	;
996	:	data_f2=	-653	;
997	:	data_f2=	-1022	;
998	:	data_f2=	-747	;
999	:	data_f2=	0	;
1000	:	data_f2=	0	;

default : data_f2=0;
endcase
always @*
case(count)
0	:	fsk_mod=	746	;
1	:	fsk_mod=	1021	;
2	:	fsk_mod=	652	;
3	:	fsk_mod=	-129	;
4	:	fsk_mod=	-829	;
5	:	fsk_mod=	-1006	;
6	:	fsk_mod=	-549	;
7	:	fsk_mod=	254	;
8	:	fsk_mod=	897	;
9	:	fsk_mod=	973	;
10	:	fsk_mod=	435	;
11	:	fsk_mod=	-377	;
12	:	fsk_mod=	-953	;
13	:	fsk_mod=	-927	;
14	:	fsk_mod=	-317	;
15	:	fsk_mod=	493	;
16	:	fsk_mod=	991	;
17	:	fsk_mod=	864	;
18	:	fsk_mod=	191	;
19	:	fsk_mod=	-602	;
20	:	fsk_mod=	-1016	;
21	:	fsk_mod=	-790	;
22	:	fsk_mod=	-65	;
23	:	fsk_mod=	700	;
24	:	fsk_mod=	1024	;
25	:	fsk_mod=	700	;
26	:	fsk_mod=	-65	;
27	:	fsk_mod=	-790	;
28	:	fsk_mod=	-1016	;
29	:	fsk_mod=	-602	;
30	:	fsk_mod=	191	;
31	:	fsk_mod=	864	;
32	:	fsk_mod=	991	;
33	:	fsk_mod=	493	;
34	:	fsk_mod=	-317	;
35	:	fsk_mod=	-927	;
36	:	fsk_mod=	-953	;
37	:	fsk_mod=	-377	;
38	:	fsk_mod=	435	;
39	:	fsk_mod=	973	;
40	:	fsk_mod=	897	;
41	:	fsk_mod=	254	;
42	:	fsk_mod=	-549	;
43	:	fsk_mod=	-1006	;
44	:	fsk_mod=	-829	;
45	:	fsk_mod=	-129	;
46	:	fsk_mod=	652	;
47	:	fsk_mod=	1021	;
48	:	fsk_mod=	746	;
49	:	fsk_mod=	-1	;
50	:	fsk_mod=	-747	;
51	:	fsk_mod=	-1022	;
52	:	fsk_mod=	-653	;
53	:	fsk_mod=	128	;
54	:	fsk_mod=	828	;
55	:	fsk_mod=	1005	;
56	:	fsk_mod=	548	;
57	:	fsk_mod=	-255	;
58	:	fsk_mod=	-898	;
59	:	fsk_mod=	-974	;
60	:	fsk_mod=	-436	;
61	:	fsk_mod=	376	;
62	:	fsk_mod=	952	;
63	:	fsk_mod=	926	;
64	:	fsk_mod=	316	;
65	:	fsk_mod=	-494	;
66	:	fsk_mod=	-992	;
67	:	fsk_mod=	-865	;
68	:	fsk_mod=	-192	;
69	:	fsk_mod=	601	;
70	:	fsk_mod=	1015	;
71	:	fsk_mod=	789	;
72	:	fsk_mod=	64	;
73	:	fsk_mod=	-701	;
74	:	fsk_mod=	-1024	;
75	:	fsk_mod=	-701	;
76	:	fsk_mod=	64	;
77	:	fsk_mod=	789	;
78	:	fsk_mod=	1015	;
79	:	fsk_mod=	601	;
80	:	fsk_mod=	-192	;
81	:	fsk_mod=	-865	;
82	:	fsk_mod=	-992	;
83	:	fsk_mod=	-494	;
84	:	fsk_mod=	316	;
85	:	fsk_mod=	926	;
86	:	fsk_mod=	952	;
87	:	fsk_mod=	376	;
88	:	fsk_mod=	-436	;
89	:	fsk_mod=	-974	;
90	:	fsk_mod=	-898	;
91	:	fsk_mod=	-255	;
92	:	fsk_mod=	548	;
93	:	fsk_mod=	1005	;
94	:	fsk_mod=	828	;
95	:	fsk_mod=	128	;
96	:	fsk_mod=	-653	;
97	:	fsk_mod=	-1022	;
98	:	fsk_mod=	-747	;
99	:	fsk_mod=	0	;
100	:	fsk_mod=	864	;
101	:	fsk_mod=	926	;
102	:	fsk_mod=	128	;
103	:	fsk_mod=	-790	;
104	:	fsk_mod=	-974	;
105	:	fsk_mod=	-255	;
106	:	fsk_mod=	700	;
107	:	fsk_mod=	1005	;
108	:	fsk_mod=	376	;
109	:	fsk_mod=	-602	;
110	:	fsk_mod=	-1022	;
111	:	fsk_mod=	-494	;
112	:	fsk_mod=	493	;
113	:	fsk_mod=	1021	;
114	:	fsk_mod=	601	;
115	:	fsk_mod=	-377	;
116	:	fsk_mod=	-1006	;
117	:	fsk_mod=	-701	;
118	:	fsk_mod=	254	;
119	:	fsk_mod=	973	;
120	:	fsk_mod=	789	;
121	:	fsk_mod=	-129	;
122	:	fsk_mod=	-927	;
123	:	fsk_mod=	-865	;
124	:	fsk_mod=	0	;
125	:	fsk_mod=	864	;
126	:	fsk_mod=	926	;
127	:	fsk_mod=	128	;
128	:	fsk_mod=	-790	;
129	:	fsk_mod=	-974	;
130	:	fsk_mod=	-255	;
131	:	fsk_mod=	700	;
132	:	fsk_mod=	1005	;
133	:	fsk_mod=	376	;
134	:	fsk_mod=	-602	;
135	:	fsk_mod=	-1022	;
136	:	fsk_mod=	-494	;
137	:	fsk_mod=	493	;
138	:	fsk_mod=	1021	;
139	:	fsk_mod=	601	;
140	:	fsk_mod=	-377	;
141	:	fsk_mod=	-1006	;
142	:	fsk_mod=	-701	;
143	:	fsk_mod=	254	;
144	:	fsk_mod=	973	;
145	:	fsk_mod=	789	;
146	:	fsk_mod=	-129	;
147	:	fsk_mod=	-927	;
148	:	fsk_mod=	-865	;
149	:	fsk_mod=	0	;
150	:	fsk_mod=	864	;
151	:	fsk_mod=	926	;
152	:	fsk_mod=	128	;
153	:	fsk_mod=	-790	;
154	:	fsk_mod=	-974	;
155	:	fsk_mod=	-255	;
156	:	fsk_mod=	700	;
157	:	fsk_mod=	1005	;
158	:	fsk_mod=	376	;
159	:	fsk_mod=	-602	;
160	:	fsk_mod=	-1022	;
161	:	fsk_mod=	-494	;
162	:	fsk_mod=	493	;
163	:	fsk_mod=	1021	;
164	:	fsk_mod=	601	;
165	:	fsk_mod=	-377	;
166	:	fsk_mod=	-1006	;
167	:	fsk_mod=	-701	;
168	:	fsk_mod=	254	;
169	:	fsk_mod=	973	;
170	:	fsk_mod=	789	;
171	:	fsk_mod=	-129	;
172	:	fsk_mod=	-927	;
173	:	fsk_mod=	-865	;
174	:	fsk_mod=	-1	;
175	:	fsk_mod=	864	;
176	:	fsk_mod=	926	;
177	:	fsk_mod=	128	;
178	:	fsk_mod=	-790	;
179	:	fsk_mod=	-974	;
180	:	fsk_mod=	-255	;
181	:	fsk_mod=	700	;
182	:	fsk_mod=	1005	;
183	:	fsk_mod=	376	;
184	:	fsk_mod=	-602	;
185	:	fsk_mod=	-1022	;
186	:	fsk_mod=	-494	;
187	:	fsk_mod=	493	;
188	:	fsk_mod=	1021	;
189	:	fsk_mod=	601	;
190	:	fsk_mod=	-377	;
191	:	fsk_mod=	-1006	;
192	:	fsk_mod=	-701	;
193	:	fsk_mod=	254	;
194	:	fsk_mod=	973	;
195	:	fsk_mod=	789	;
196	:	fsk_mod=	-129	;
197	:	fsk_mod=	-927	;
198	:	fsk_mod=	-865	;
199	:	fsk_mod=	-1	;
200	:	fsk_mod=	746	;
201	:	fsk_mod=	1021	;
202	:	fsk_mod=	652	;
203	:	fsk_mod=	-129	;
204	:	fsk_mod=	-829	;
205	:	fsk_mod=	-1006	;
206	:	fsk_mod=	-549	;
207	:	fsk_mod=	254	;
208	:	fsk_mod=	897	;
209	:	fsk_mod=	973	;
210	:	fsk_mod=	435	;
211	:	fsk_mod=	-377	;
212	:	fsk_mod=	-953	;
213	:	fsk_mod=	-927	;
214	:	fsk_mod=	-317	;
215	:	fsk_mod=	493	;
216	:	fsk_mod=	991	;
217	:	fsk_mod=	864	;
218	:	fsk_mod=	191	;
219	:	fsk_mod=	-602	;
220	:	fsk_mod=	-1016	;
221	:	fsk_mod=	-790	;
222	:	fsk_mod=	-65	;
223	:	fsk_mod=	700	;
224	:	fsk_mod=	1024	;
225	:	fsk_mod=	700	;
226	:	fsk_mod=	-65	;
227	:	fsk_mod=	-790	;
228	:	fsk_mod=	-1016	;
229	:	fsk_mod=	-602	;
230	:	fsk_mod=	191	;
231	:	fsk_mod=	864	;
232	:	fsk_mod=	991	;
233	:	fsk_mod=	493	;
234	:	fsk_mod=	-317	;
235	:	fsk_mod=	-927	;
236	:	fsk_mod=	-953	;
237	:	fsk_mod=	-377	;
238	:	fsk_mod=	435	;
239	:	fsk_mod=	973	;
240	:	fsk_mod=	897	;
241	:	fsk_mod=	254	;
242	:	fsk_mod=	-549	;
243	:	fsk_mod=	-1006	;
244	:	fsk_mod=	-829	;
245	:	fsk_mod=	-129	;
246	:	fsk_mod=	652	;
247	:	fsk_mod=	1021	;
248	:	fsk_mod=	746	;
249	:	fsk_mod=	-1	;
250	:	fsk_mod=	-747	;
251	:	fsk_mod=	-1022	;
252	:	fsk_mod=	-653	;
253	:	fsk_mod=	128	;
254	:	fsk_mod=	828	;
255	:	fsk_mod=	1005	;
256	:	fsk_mod=	548	;
257	:	fsk_mod=	-255	;
258	:	fsk_mod=	-898	;
259	:	fsk_mod=	-974	;
260	:	fsk_mod=	-436	;
261	:	fsk_mod=	376	;
262	:	fsk_mod=	952	;
263	:	fsk_mod=	926	;
264	:	fsk_mod=	316	;
265	:	fsk_mod=	-494	;
266	:	fsk_mod=	-992	;
267	:	fsk_mod=	-865	;
268	:	fsk_mod=	-192	;
269	:	fsk_mod=	601	;
270	:	fsk_mod=	1015	;
271	:	fsk_mod=	789	;
272	:	fsk_mod=	64	;
273	:	fsk_mod=	-701	;
274	:	fsk_mod=	-1024	;
275	:	fsk_mod=	-701	;
276	:	fsk_mod=	64	;
277	:	fsk_mod=	789	;
278	:	fsk_mod=	1015	;
279	:	fsk_mod=	601	;
280	:	fsk_mod=	-192	;
281	:	fsk_mod=	-865	;
282	:	fsk_mod=	-992	;
283	:	fsk_mod=	-494	;
284	:	fsk_mod=	316	;
285	:	fsk_mod=	926	;
286	:	fsk_mod=	952	;
287	:	fsk_mod=	376	;
288	:	fsk_mod=	-436	;
289	:	fsk_mod=	-974	;
290	:	fsk_mod=	-898	;
291	:	fsk_mod=	-255	;
292	:	fsk_mod=	548	;
293	:	fsk_mod=	1005	;
294	:	fsk_mod=	828	;
295	:	fsk_mod=	128	;
296	:	fsk_mod=	-653	;
297	:	fsk_mod=	-1022	;
298	:	fsk_mod=	-747	;
299	:	fsk_mod=	0	;
300	:	fsk_mod=	746	;
301	:	fsk_mod=	1021	;
302	:	fsk_mod=	652	;
303	:	fsk_mod=	-129	;
304	:	fsk_mod=	-829	;
305	:	fsk_mod=	-1006	;
306	:	fsk_mod=	-549	;
307	:	fsk_mod=	254	;
308	:	fsk_mod=	897	;
309	:	fsk_mod=	973	;
310	:	fsk_mod=	435	;
311	:	fsk_mod=	-377	;
312	:	fsk_mod=	-953	;
313	:	fsk_mod=	-927	;
314	:	fsk_mod=	-317	;
315	:	fsk_mod=	493	;
316	:	fsk_mod=	991	;
317	:	fsk_mod=	864	;
318	:	fsk_mod=	191	;
319	:	fsk_mod=	-602	;
320	:	fsk_mod=	-1016	;
321	:	fsk_mod=	-790	;
322	:	fsk_mod=	-65	;
323	:	fsk_mod=	700	;
324	:	fsk_mod=	1024	;
325	:	fsk_mod=	700	;
326	:	fsk_mod=	-65	;
327	:	fsk_mod=	-790	;
328	:	fsk_mod=	-1016	;
329	:	fsk_mod=	-602	;
330	:	fsk_mod=	191	;
331	:	fsk_mod=	864	;
332	:	fsk_mod=	991	;
333	:	fsk_mod=	493	;
334	:	fsk_mod=	-317	;
335	:	fsk_mod=	-927	;
336	:	fsk_mod=	-953	;
337	:	fsk_mod=	-377	;
338	:	fsk_mod=	435	;
339	:	fsk_mod=	973	;
340	:	fsk_mod=	897	;
341	:	fsk_mod=	254	;
342	:	fsk_mod=	-549	;
343	:	fsk_mod=	-1006	;
344	:	fsk_mod=	-829	;
345	:	fsk_mod=	-129	;
346	:	fsk_mod=	652	;
347	:	fsk_mod=	1021	;
348	:	fsk_mod=	746	;
349	:	fsk_mod=	-1	;
350	:	fsk_mod=	-747	;
351	:	fsk_mod=	-1022	;
352	:	fsk_mod=	-653	;
353	:	fsk_mod=	128	;
354	:	fsk_mod=	828	;
355	:	fsk_mod=	1005	;
356	:	fsk_mod=	548	;
357	:	fsk_mod=	-255	;
358	:	fsk_mod=	-898	;
359	:	fsk_mod=	-974	;
360	:	fsk_mod=	-436	;
361	:	fsk_mod=	376	;
362	:	fsk_mod=	952	;
363	:	fsk_mod=	926	;
364	:	fsk_mod=	316	;
365	:	fsk_mod=	-494	;
366	:	fsk_mod=	-992	;
367	:	fsk_mod=	-865	;
368	:	fsk_mod=	-192	;
369	:	fsk_mod=	601	;
370	:	fsk_mod=	1015	;
371	:	fsk_mod=	789	;
372	:	fsk_mod=	64	;
373	:	fsk_mod=	-701	;
374	:	fsk_mod=	-1024	;
375	:	fsk_mod=	-701	;
376	:	fsk_mod=	64	;
377	:	fsk_mod=	789	;
378	:	fsk_mod=	1015	;
379	:	fsk_mod=	601	;
380	:	fsk_mod=	-192	;
381	:	fsk_mod=	-865	;
382	:	fsk_mod=	-992	;
383	:	fsk_mod=	-494	;
384	:	fsk_mod=	316	;
385	:	fsk_mod=	926	;
386	:	fsk_mod=	952	;
387	:	fsk_mod=	376	;
388	:	fsk_mod=	-436	;
389	:	fsk_mod=	-974	;
390	:	fsk_mod=	-898	;
391	:	fsk_mod=	-255	;
392	:	fsk_mod=	548	;
393	:	fsk_mod=	1005	;
394	:	fsk_mod=	828	;
395	:	fsk_mod=	128	;
396	:	fsk_mod=	-653	;
397	:	fsk_mod=	-1022	;
398	:	fsk_mod=	-747	;
399	:	fsk_mod=	0	;
400	:	fsk_mod=	864	;
401	:	fsk_mod=	926	;
402	:	fsk_mod=	128	;
403	:	fsk_mod=	-790	;
404	:	fsk_mod=	-974	;
405	:	fsk_mod=	-255	;
406	:	fsk_mod=	700	;
407	:	fsk_mod=	1005	;
408	:	fsk_mod=	376	;
409	:	fsk_mod=	-602	;
410	:	fsk_mod=	-1022	;
411	:	fsk_mod=	-494	;
412	:	fsk_mod=	493	;
413	:	fsk_mod=	1021	;
414	:	fsk_mod=	601	;
415	:	fsk_mod=	-377	;
416	:	fsk_mod=	-1006	;
417	:	fsk_mod=	-701	;
418	:	fsk_mod=	254	;
419	:	fsk_mod=	973	;
420	:	fsk_mod=	789	;
421	:	fsk_mod=	-129	;
422	:	fsk_mod=	-927	;
423	:	fsk_mod=	-865	;
424	:	fsk_mod=	0	;
425	:	fsk_mod=	864	;
426	:	fsk_mod=	926	;
427	:	fsk_mod=	128	;
428	:	fsk_mod=	-790	;
429	:	fsk_mod=	-974	;
430	:	fsk_mod=	-255	;
431	:	fsk_mod=	700	;
432	:	fsk_mod=	1005	;
433	:	fsk_mod=	376	;
434	:	fsk_mod=	-602	;
435	:	fsk_mod=	-1022	;
436	:	fsk_mod=	-494	;
437	:	fsk_mod=	493	;
438	:	fsk_mod=	1021	;
439	:	fsk_mod=	601	;
440	:	fsk_mod=	-377	;
441	:	fsk_mod=	-1006	;
442	:	fsk_mod=	-701	;
443	:	fsk_mod=	254	;
444	:	fsk_mod=	973	;
445	:	fsk_mod=	789	;
446	:	fsk_mod=	-129	;
447	:	fsk_mod=	-927	;
448	:	fsk_mod=	-865	;
449	:	fsk_mod=	0	;
450	:	fsk_mod=	864	;
451	:	fsk_mod=	926	;
452	:	fsk_mod=	128	;
453	:	fsk_mod=	-790	;
454	:	fsk_mod=	-974	;
455	:	fsk_mod=	-255	;
456	:	fsk_mod=	700	;
457	:	fsk_mod=	1005	;
458	:	fsk_mod=	376	;
459	:	fsk_mod=	-602	;
460	:	fsk_mod=	-1022	;
461	:	fsk_mod=	-494	;
462	:	fsk_mod=	493	;
463	:	fsk_mod=	1021	;
464	:	fsk_mod=	601	;
465	:	fsk_mod=	-377	;
466	:	fsk_mod=	-1006	;
467	:	fsk_mod=	-701	;
468	:	fsk_mod=	254	;
469	:	fsk_mod=	973	;
470	:	fsk_mod=	789	;
471	:	fsk_mod=	-129	;
472	:	fsk_mod=	-927	;
473	:	fsk_mod=	-865	;
474	:	fsk_mod=	-1	;
475	:	fsk_mod=	864	;
476	:	fsk_mod=	926	;
477	:	fsk_mod=	128	;
478	:	fsk_mod=	-790	;
479	:	fsk_mod=	-974	;
480	:	fsk_mod=	-255	;
481	:	fsk_mod=	700	;
482	:	fsk_mod=	1005	;
483	:	fsk_mod=	376	;
484	:	fsk_mod=	-602	;
485	:	fsk_mod=	-1022	;
486	:	fsk_mod=	-494	;
487	:	fsk_mod=	493	;
488	:	fsk_mod=	1021	;
489	:	fsk_mod=	601	;
490	:	fsk_mod=	-377	;
491	:	fsk_mod=	-1006	;
492	:	fsk_mod=	-701	;
493	:	fsk_mod=	254	;
494	:	fsk_mod=	973	;
495	:	fsk_mod=	789	;
496	:	fsk_mod=	-129	;
497	:	fsk_mod=	-927	;
498	:	fsk_mod=	-865	;
499	:	fsk_mod=	-1	;
500	:	fsk_mod=	746	;
501	:	fsk_mod=	1021	;
502	:	fsk_mod=	652	;
503	:	fsk_mod=	-129	;
504	:	fsk_mod=	-829	;
505	:	fsk_mod=	-1006	;
506	:	fsk_mod=	-549	;
507	:	fsk_mod=	254	;
508	:	fsk_mod=	897	;
509	:	fsk_mod=	973	;
510	:	fsk_mod=	435	;
511	:	fsk_mod=	-377	;
512	:	fsk_mod=	-953	;
513	:	fsk_mod=	-927	;
514	:	fsk_mod=	-317	;
515	:	fsk_mod=	493	;
516	:	fsk_mod=	991	;
517	:	fsk_mod=	864	;
518	:	fsk_mod=	191	;
519	:	fsk_mod=	-602	;
520	:	fsk_mod=	-1016	;
521	:	fsk_mod=	-790	;
522	:	fsk_mod=	-65	;
523	:	fsk_mod=	700	;
524	:	fsk_mod=	1024	;
525	:	fsk_mod=	700	;
526	:	fsk_mod=	-65	;
527	:	fsk_mod=	-790	;
528	:	fsk_mod=	-1016	;
529	:	fsk_mod=	-602	;
530	:	fsk_mod=	191	;
531	:	fsk_mod=	864	;
532	:	fsk_mod=	991	;
533	:	fsk_mod=	493	;
534	:	fsk_mod=	-317	;
535	:	fsk_mod=	-927	;
536	:	fsk_mod=	-953	;
537	:	fsk_mod=	-377	;
538	:	fsk_mod=	435	;
539	:	fsk_mod=	973	;
540	:	fsk_mod=	897	;
541	:	fsk_mod=	254	;
542	:	fsk_mod=	-549	;
543	:	fsk_mod=	-1006	;
544	:	fsk_mod=	-829	;
545	:	fsk_mod=	-129	;
546	:	fsk_mod=	652	;
547	:	fsk_mod=	1021	;
548	:	fsk_mod=	746	;
549	:	fsk_mod=	-1	;
550	:	fsk_mod=	-747	;
551	:	fsk_mod=	-1022	;
552	:	fsk_mod=	-653	;
553	:	fsk_mod=	128	;
554	:	fsk_mod=	828	;
555	:	fsk_mod=	1005	;
556	:	fsk_mod=	548	;
557	:	fsk_mod=	-255	;
558	:	fsk_mod=	-898	;
559	:	fsk_mod=	-974	;
560	:	fsk_mod=	-436	;
561	:	fsk_mod=	376	;
562	:	fsk_mod=	952	;
563	:	fsk_mod=	926	;
564	:	fsk_mod=	316	;
565	:	fsk_mod=	-494	;
566	:	fsk_mod=	-992	;
567	:	fsk_mod=	-865	;
568	:	fsk_mod=	-192	;
569	:	fsk_mod=	601	;
570	:	fsk_mod=	1015	;
571	:	fsk_mod=	789	;
572	:	fsk_mod=	64	;
573	:	fsk_mod=	-701	;
574	:	fsk_mod=	-1024	;
575	:	fsk_mod=	-701	;
576	:	fsk_mod=	64	;
577	:	fsk_mod=	789	;
578	:	fsk_mod=	1015	;
579	:	fsk_mod=	601	;
580	:	fsk_mod=	-192	;
581	:	fsk_mod=	-865	;
582	:	fsk_mod=	-992	;
583	:	fsk_mod=	-494	;
584	:	fsk_mod=	316	;
585	:	fsk_mod=	926	;
586	:	fsk_mod=	952	;
587	:	fsk_mod=	376	;
588	:	fsk_mod=	-436	;
589	:	fsk_mod=	-974	;
590	:	fsk_mod=	-898	;
591	:	fsk_mod=	-255	;
592	:	fsk_mod=	548	;
593	:	fsk_mod=	1005	;
594	:	fsk_mod=	828	;
595	:	fsk_mod=	128	;
596	:	fsk_mod=	-653	;
597	:	fsk_mod=	-1022	;
598	:	fsk_mod=	-747	;
599	:	fsk_mod=	0	;
600	:	fsk_mod=	864	;
601	:	fsk_mod=	926	;
602	:	fsk_mod=	128	;
603	:	fsk_mod=	-790	;
604	:	fsk_mod=	-974	;
605	:	fsk_mod=	-255	;
606	:	fsk_mod=	700	;
607	:	fsk_mod=	1005	;
608	:	fsk_mod=	376	;
609	:	fsk_mod=	-602	;
610	:	fsk_mod=	-1022	;
611	:	fsk_mod=	-494	;
612	:	fsk_mod=	493	;
613	:	fsk_mod=	1021	;
614	:	fsk_mod=	601	;
615	:	fsk_mod=	-377	;
616	:	fsk_mod=	-1006	;
617	:	fsk_mod=	-701	;
618	:	fsk_mod=	254	;
619	:	fsk_mod=	973	;
620	:	fsk_mod=	789	;
621	:	fsk_mod=	-129	;
622	:	fsk_mod=	-927	;
623	:	fsk_mod=	-865	;
624	:	fsk_mod=	0	;
625	:	fsk_mod=	864	;
626	:	fsk_mod=	926	;
627	:	fsk_mod=	128	;
628	:	fsk_mod=	-790	;
629	:	fsk_mod=	-974	;
630	:	fsk_mod=	-255	;
631	:	fsk_mod=	700	;
632	:	fsk_mod=	1005	;
633	:	fsk_mod=	376	;
634	:	fsk_mod=	-602	;
635	:	fsk_mod=	-1022	;
636	:	fsk_mod=	-494	;
637	:	fsk_mod=	493	;
638	:	fsk_mod=	1021	;
639	:	fsk_mod=	601	;
640	:	fsk_mod=	-377	;
641	:	fsk_mod=	-1006	;
642	:	fsk_mod=	-701	;
643	:	fsk_mod=	254	;
644	:	fsk_mod=	973	;
645	:	fsk_mod=	789	;
646	:	fsk_mod=	-129	;
647	:	fsk_mod=	-927	;
648	:	fsk_mod=	-865	;
649	:	fsk_mod=	0	;
650	:	fsk_mod=	864	;
651	:	fsk_mod=	926	;
652	:	fsk_mod=	128	;
653	:	fsk_mod=	-790	;
654	:	fsk_mod=	-974	;
655	:	fsk_mod=	-255	;
656	:	fsk_mod=	700	;
657	:	fsk_mod=	1005	;
658	:	fsk_mod=	376	;
659	:	fsk_mod=	-602	;
660	:	fsk_mod=	-1022	;
661	:	fsk_mod=	-494	;
662	:	fsk_mod=	493	;
663	:	fsk_mod=	1021	;
664	:	fsk_mod=	601	;
665	:	fsk_mod=	-377	;
666	:	fsk_mod=	-1006	;
667	:	fsk_mod=	-701	;
668	:	fsk_mod=	254	;
669	:	fsk_mod=	973	;
670	:	fsk_mod=	789	;
671	:	fsk_mod=	-129	;
672	:	fsk_mod=	-927	;
673	:	fsk_mod=	-865	;
674	:	fsk_mod=	-1	;
675	:	fsk_mod=	864	;
676	:	fsk_mod=	926	;
677	:	fsk_mod=	128	;
678	:	fsk_mod=	-790	;
679	:	fsk_mod=	-974	;
680	:	fsk_mod=	-255	;
681	:	fsk_mod=	700	;
682	:	fsk_mod=	1005	;
683	:	fsk_mod=	376	;
684	:	fsk_mod=	-602	;
685	:	fsk_mod=	-1022	;
686	:	fsk_mod=	-494	;
687	:	fsk_mod=	493	;
688	:	fsk_mod=	1021	;
689	:	fsk_mod=	601	;
690	:	fsk_mod=	-377	;
691	:	fsk_mod=	-1006	;
692	:	fsk_mod=	-701	;
693	:	fsk_mod=	254	;
694	:	fsk_mod=	973	;
695	:	fsk_mod=	789	;
696	:	fsk_mod=	-129	;
697	:	fsk_mod=	-927	;
698	:	fsk_mod=	-865	;
699	:	fsk_mod=	-1	;
700	:	fsk_mod=	864	;
701	:	fsk_mod=	926	;
702	:	fsk_mod=	128	;
703	:	fsk_mod=	-790	;
704	:	fsk_mod=	-974	;
705	:	fsk_mod=	-255	;
706	:	fsk_mod=	700	;
707	:	fsk_mod=	1005	;
708	:	fsk_mod=	376	;
709	:	fsk_mod=	-602	;
710	:	fsk_mod=	-1022	;
711	:	fsk_mod=	-494	;
712	:	fsk_mod=	493	;
713	:	fsk_mod=	1021	;
714	:	fsk_mod=	601	;
715	:	fsk_mod=	-377	;
716	:	fsk_mod=	-1006	;
717	:	fsk_mod=	-701	;
718	:	fsk_mod=	254	;
719	:	fsk_mod=	973	;
720	:	fsk_mod=	789	;
721	:	fsk_mod=	-129	;
722	:	fsk_mod=	-927	;
723	:	fsk_mod=	-865	;
724	:	fsk_mod=	0	;
725	:	fsk_mod=	864	;
726	:	fsk_mod=	926	;
727	:	fsk_mod=	128	;
728	:	fsk_mod=	-790	;
729	:	fsk_mod=	-974	;
730	:	fsk_mod=	-255	;
731	:	fsk_mod=	700	;
732	:	fsk_mod=	1005	;
733	:	fsk_mod=	376	;
734	:	fsk_mod=	-602	;
735	:	fsk_mod=	-1022	;
736	:	fsk_mod=	-494	;
737	:	fsk_mod=	493	;
738	:	fsk_mod=	1021	;
739	:	fsk_mod=	601	;
740	:	fsk_mod=	-377	;
741	:	fsk_mod=	-1006	;
742	:	fsk_mod=	-701	;
743	:	fsk_mod=	254	;
744	:	fsk_mod=	973	;
745	:	fsk_mod=	789	;
746	:	fsk_mod=	-129	;
747	:	fsk_mod=	-927	;
748	:	fsk_mod=	-865	;
749	:	fsk_mod=	0	;
750	:	fsk_mod=	864	;
751	:	fsk_mod=	926	;
752	:	fsk_mod=	128	;
753	:	fsk_mod=	-790	;
754	:	fsk_mod=	-974	;
755	:	fsk_mod=	-255	;
756	:	fsk_mod=	700	;
757	:	fsk_mod=	1005	;
758	:	fsk_mod=	376	;
759	:	fsk_mod=	-602	;
760	:	fsk_mod=	-1022	;
761	:	fsk_mod=	-494	;
762	:	fsk_mod=	493	;
763	:	fsk_mod=	1021	;
764	:	fsk_mod=	601	;
765	:	fsk_mod=	-377	;
766	:	fsk_mod=	-1006	;
767	:	fsk_mod=	-701	;
768	:	fsk_mod=	254	;
769	:	fsk_mod=	973	;
770	:	fsk_mod=	789	;
771	:	fsk_mod=	-129	;
772	:	fsk_mod=	-927	;
773	:	fsk_mod=	-865	;
774	:	fsk_mod=	-1	;
775	:	fsk_mod=	864	;
776	:	fsk_mod=	926	;
777	:	fsk_mod=	128	;
778	:	fsk_mod=	-790	;
779	:	fsk_mod=	-974	;
780	:	fsk_mod=	-255	;
781	:	fsk_mod=	700	;
782	:	fsk_mod=	1005	;
783	:	fsk_mod=	376	;
784	:	fsk_mod=	-602	;
785	:	fsk_mod=	-1022	;
786	:	fsk_mod=	-494	;
787	:	fsk_mod=	493	;
788	:	fsk_mod=	1021	;
789	:	fsk_mod=	601	;
790	:	fsk_mod=	-377	;
791	:	fsk_mod=	-1006	;
792	:	fsk_mod=	-701	;
793	:	fsk_mod=	254	;
794	:	fsk_mod=	973	;
795	:	fsk_mod=	789	;
796	:	fsk_mod=	-129	;
797	:	fsk_mod=	-927	;
798	:	fsk_mod=	-865	;
799	:	fsk_mod=	-1	;
800	:	fsk_mod=	746	;
801	:	fsk_mod=	1021	;
802	:	fsk_mod=	652	;
803	:	fsk_mod=	-129	;
804	:	fsk_mod=	-829	;
805	:	fsk_mod=	-1006	;
806	:	fsk_mod=	-549	;
807	:	fsk_mod=	254	;
808	:	fsk_mod=	897	;
809	:	fsk_mod=	973	;
810	:	fsk_mod=	435	;
811	:	fsk_mod=	-377	;
812	:	fsk_mod=	-953	;
813	:	fsk_mod=	-927	;
814	:	fsk_mod=	-317	;
815	:	fsk_mod=	493	;
816	:	fsk_mod=	991	;
817	:	fsk_mod=	864	;
818	:	fsk_mod=	191	;
819	:	fsk_mod=	-602	;
820	:	fsk_mod=	-1016	;
821	:	fsk_mod=	-790	;
822	:	fsk_mod=	-65	;
823	:	fsk_mod=	700	;
824	:	fsk_mod=	1024	;
825	:	fsk_mod=	700	;
826	:	fsk_mod=	-65	;
827	:	fsk_mod=	-790	;
828	:	fsk_mod=	-1016	;
829	:	fsk_mod=	-602	;
830	:	fsk_mod=	191	;
831	:	fsk_mod=	864	;
832	:	fsk_mod=	991	;
833	:	fsk_mod=	493	;
834	:	fsk_mod=	-317	;
835	:	fsk_mod=	-927	;
836	:	fsk_mod=	-953	;
837	:	fsk_mod=	-377	;
838	:	fsk_mod=	435	;
839	:	fsk_mod=	973	;
840	:	fsk_mod=	897	;
841	:	fsk_mod=	254	;
842	:	fsk_mod=	-549	;
843	:	fsk_mod=	-1006	;
844	:	fsk_mod=	-829	;
845	:	fsk_mod=	-129	;
846	:	fsk_mod=	652	;
847	:	fsk_mod=	1021	;
848	:	fsk_mod=	746	;
849	:	fsk_mod=	-1	;
850	:	fsk_mod=	-747	;
851	:	fsk_mod=	-1022	;
852	:	fsk_mod=	-653	;
853	:	fsk_mod=	128	;
854	:	fsk_mod=	828	;
855	:	fsk_mod=	1005	;
856	:	fsk_mod=	548	;
857	:	fsk_mod=	-255	;
858	:	fsk_mod=	-898	;
859	:	fsk_mod=	-974	;
860	:	fsk_mod=	-436	;
861	:	fsk_mod=	376	;
862	:	fsk_mod=	952	;
863	:	fsk_mod=	926	;
864	:	fsk_mod=	316	;
865	:	fsk_mod=	-494	;
866	:	fsk_mod=	-992	;
867	:	fsk_mod=	-865	;
868	:	fsk_mod=	-192	;
869	:	fsk_mod=	601	;
870	:	fsk_mod=	1015	;
871	:	fsk_mod=	789	;
872	:	fsk_mod=	64	;
873	:	fsk_mod=	-701	;
874	:	fsk_mod=	-1024	;
875	:	fsk_mod=	-701	;
876	:	fsk_mod=	64	;
877	:	fsk_mod=	789	;
878	:	fsk_mod=	1015	;
879	:	fsk_mod=	601	;
880	:	fsk_mod=	-192	;
881	:	fsk_mod=	-865	;
882	:	fsk_mod=	-992	;
883	:	fsk_mod=	-494	;
884	:	fsk_mod=	316	;
885	:	fsk_mod=	926	;
886	:	fsk_mod=	952	;
887	:	fsk_mod=	376	;
888	:	fsk_mod=	-436	;
889	:	fsk_mod=	-974	;
890	:	fsk_mod=	-898	;
891	:	fsk_mod=	-255	;
892	:	fsk_mod=	548	;
893	:	fsk_mod=	1005	;
894	:	fsk_mod=	828	;
895	:	fsk_mod=	128	;
896	:	fsk_mod=	-653	;
897	:	fsk_mod=	-1022	;
898	:	fsk_mod=	-747	;
899	:	fsk_mod=	0	;
900	:	fsk_mod=	746	;
901	:	fsk_mod=	1021	;
902	:	fsk_mod=	652	;
903	:	fsk_mod=	-129	;
904	:	fsk_mod=	-829	;
905	:	fsk_mod=	-1006	;
906	:	fsk_mod=	-549	;
907	:	fsk_mod=	254	;
908	:	fsk_mod=	897	;
909	:	fsk_mod=	973	;
910	:	fsk_mod=	435	;
911	:	fsk_mod=	-377	;
912	:	fsk_mod=	-953	;
913	:	fsk_mod=	-927	;
914	:	fsk_mod=	-317	;
915	:	fsk_mod=	493	;
916	:	fsk_mod=	991	;
917	:	fsk_mod=	864	;
918	:	fsk_mod=	191	;
919	:	fsk_mod=	-602	;
920	:	fsk_mod=	-1016	;
921	:	fsk_mod=	-790	;
922	:	fsk_mod=	-65	;
923	:	fsk_mod=	700	;
924	:	fsk_mod=	1024	;
925	:	fsk_mod=	700	;
926	:	fsk_mod=	-65	;
927	:	fsk_mod=	-790	;
928	:	fsk_mod=	-1016	;
929	:	fsk_mod=	-602	;
930	:	fsk_mod=	191	;
931	:	fsk_mod=	864	;
932	:	fsk_mod=	991	;
933	:	fsk_mod=	493	;
934	:	fsk_mod=	-317	;
935	:	fsk_mod=	-927	;
936	:	fsk_mod=	-953	;
937	:	fsk_mod=	-377	;
938	:	fsk_mod=	435	;
939	:	fsk_mod=	973	;
940	:	fsk_mod=	897	;
941	:	fsk_mod=	254	;
942	:	fsk_mod=	-549	;
943	:	fsk_mod=	-1006	;
944	:	fsk_mod=	-829	;
945	:	fsk_mod=	-129	;
946	:	fsk_mod=	652	;
947	:	fsk_mod=	1021	;
948	:	fsk_mod=	746	;
949	:	fsk_mod=	-1	;
950	:	fsk_mod=	-747	;
951	:	fsk_mod=	-1022	;
952	:	fsk_mod=	-653	;
953	:	fsk_mod=	128	;
954	:	fsk_mod=	828	;
955	:	fsk_mod=	1005	;
956	:	fsk_mod=	548	;
957	:	fsk_mod=	-255	;
958	:	fsk_mod=	-898	;
959	:	fsk_mod=	-974	;
960	:	fsk_mod=	-436	;
961	:	fsk_mod=	376	;
962	:	fsk_mod=	952	;
963	:	fsk_mod=	926	;
964	:	fsk_mod=	316	;
965	:	fsk_mod=	-494	;
966	:	fsk_mod=	-992	;
967	:	fsk_mod=	-865	;
968	:	fsk_mod=	-192	;
969	:	fsk_mod=	601	;
970	:	fsk_mod=	1015	;
971	:	fsk_mod=	789	;
972	:	fsk_mod=	64	;
973	:	fsk_mod=	-701	;
974	:	fsk_mod=	-1024	;
975	:	fsk_mod=	-701	;
976	:	fsk_mod=	64	;
977	:	fsk_mod=	789	;
978	:	fsk_mod=	1015	;
979	:	fsk_mod=	601	;
980	:	fsk_mod=	-192	;
981	:	fsk_mod=	-865	;
982	:	fsk_mod=	-992	;
983	:	fsk_mod=	-494	;
984	:	fsk_mod=	316	;
985	:	fsk_mod=	926	;
986	:	fsk_mod=	952	;
987	:	fsk_mod=	376	;
988	:	fsk_mod=	-436	;
989	:	fsk_mod=	-974	;
990	:	fsk_mod=	-898	;
991	:	fsk_mod=	-255	;
992	:	fsk_mod=	548	;
993	:	fsk_mod=	1005	;
994	:	fsk_mod=	828	;
995	:	fsk_mod=	128	;
996	:	fsk_mod=	-653	;
997	:	fsk_mod=	-1022	;
998	:	fsk_mod=	-747	;
999	:	fsk_mod=	0	;
default : fsk_mod=0;
endcase
nhan_co_dau_16bit mul_f1(
    .a(data_f1),
    .b(fsk_mod),
    .result(temp_f1)
);
nhan_co_dau_16bit mul_f2(
    .a(data_f2),
    .b(fsk_mod),
    .result(temp_f2)
);
assign mul_signal_f1=temp_f1[25:10];
assign mul_signal_f2=temp_f2[25:10];
endmodule