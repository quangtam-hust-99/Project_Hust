module tb_demodulation;
reg clk,reset;
wire  fsk_demod;
demodulation uut(
    .clk(clk),
    .reset(reset),
    .fsk_demod(fsk_demod)
);
initial begin
  clk=1;
  reset=1;
  #20 reset=0;
end

always begin
  #5 clk=~clk;
  end
 /*			
	data_f1=	737	
	data_f2=	622	;
#8000	data_f1=	1023	
	data_f2=	988	;
#8000	data_f1=	681	
	data_f2=	947	;
#8000	data_f1=	-78	
	data_f2=	515	;
#8000	data_f1=	-790	
	data_f2=	-129	;
#8000	data_f1=	-1018	
	data_f2=	-720	;
#8000	data_f1=	-623	
	data_f2=	-1015	;
#8000	data_f1=	153	
	data_f2=	-892	;
#8000	data_f1=	835	
	data_f2=	-401	;
#8000	data_f1=	1005	
	data_f2=	254	;
#8000	data_f1=	559	
	data_f2=	805	;
#8000	data_f1=	-230	
	data_f2=	1023	;
#8000	data_f1=	-879	
	data_f2=	820	;
#8000	data_f1=	-989	
	data_f2=	279	;
#8000	data_f1=	-494	
	data_f2=	-377	;
#8000	data_f1=	304	
	data_f2=	-879	;
#8000	data_f1=	915	
	data_f2=	-1018	;
#8000	data_f1=	965	
	data_f2=	-738	;
#8000	data_f1=	424	
	data_f2=	-154	;
#8000	data_f1=	-377	
	data_f2=	493	;
#8000	data_f1=	-948	
	data_f2=	937	;
#8000	data_f1=	-938	
	data_f2=	994	;
#8000	data_f1=	-353	
	data_f2=	642	;
#8000	data_f1=	447	
	data_f2=	25	;
#8000	data_f1=	973	
	data_f2=	-602	;
#8000	data_f1=	903	
	data_f2=	-982	;
#8000	data_f1=	279	
	data_f2=	-957	;
#8000	data_f1=	-516	
	data_f2=	-538	;
#8000	data_f1=	-995	
	data_f2=	102	;
#8000	data_f1=	-865	
	data_f2=	700	;
#8000	data_f1=	-205	
	data_f2=	1010	;
#8000	data_f1=	580	
	data_f2=	903	;
#8000	data_f1=	1010	
	data_f2=	424	;
#8000	data_f1=	820	
	data_f2=	-230	;
#8000	data_f1=	128	
	data_f2=	-790	;
#8000	data_f1=	-643	
	data_f2=	-1024	;
#8000	data_f1=	-1021	
	data_f2=	-836	;
#8000	data_f1=	-773	
	data_f2=	-305	;
#8000	data_f1=	-52	
	data_f2=	352	;
#8000	data_f1=	700	
	data_f2=	864	;
#8000	data_f1=	1023	
	data_f2=	1020	;
#8000	data_f1=	719	
	data_f2=	755	;
#8000	data_f1=	-26	
	data_f2=	179	;
#8000	data_f1=	-756	
	data_f2=	-471	;
#8000	data_f1=	-1022	
	data_f2=	-927	;
#8000	data_f1=	-663	
	data_f2=	-1001	;
#8000	data_f1=	102	
	data_f2=	-663	;
#8000	data_f1=	805	
	data_f2=	-52	;
#8000	data_f1=	1014	
	data_f2=	580	;
#8000	data_f1=	601	
	data_f2=	973	;
#8000	data_f1=	-180	
	data_f2=	965	;
#8000	data_f1=	-851	
	data_f2=	559	;
#8000	data_f1=	-1001	
	data_f2=	-78	;
#8000	data_f1=	-538	
	data_f2=	-682	;
#8000	data_f1=	254	
	data_f2=	-1006	;
#8000	data_f1=	891	
	data_f2=	-916	;
#8000	data_f1=	981	
	data_f2=	-448	;
#8000	data_f1=	470	
	data_f2=	204	;
#8000	data_f1=	-329	
	data_f2=	772	;
#8000	data_f1=	-927	
	data_f2=	1021	;
#8000	data_f1=	-957	
	data_f2=	850	;
#8000	data_f1=	-401	
	data_f2=	328	;
#8000	data_f1=	400	
	data_f2=	-329	;
#8000	data_f1=	956	
	data_f2=	-850	;
#8000	data_f1=	926	
	data_f2=	-1022	;
#8000	data_f1=	328	
	data_f2=	-772	;
#8000	data_f1=	-471	
	data_f2=	-204	;
#8000	data_f1=	-982	
	data_f2=	448	;
#8000	data_f1=	-892	
	data_f2=	915	;
#8000	data_f1=	-255	
	data_f2=	1006	;
#8000	data_f1=	537	
	data_f2=	682	;
#8000	data_f1=	1000	
	data_f2=	77	;
#8000	data_f1=	850	
	data_f2=	-560	;
#8000	data_f1=	179	
	data_f2=	-965	;
#8000	data_f1=	-602	
	data_f2=	-974	;
#8000	data_f1=	-1015	
	data_f2=	-581	;
#8000	data_f1=	-806	
	data_f2=	51	;
#8000	data_f1=	-103	
	data_f2=	663	;
#8000	data_f1=	662	
	data_f2=	1001	;
#8000	data_f1=	1021	
	data_f2=	926	;
#8000	data_f1=	755	
	data_f2=	471	;
#8000	data_f1=	25	
	data_f2=	-179	;
#8000	data_f1=	-720	
	data_f2=	-755	;
#8000	data_f1=	-1024	
	data_f2=	-1020	;
#8000	data_f1=	-701	
	data_f2=	-864	;
#8000	data_f1=	51	
	data_f2=	-352	;
#8000	data_f1=	772	
	data_f2=	304	;
#8000	data_f1=	1020	
	data_f2=	836	;
#8000	data_f1=	642	
	data_f2=	1023	;
#8000	data_f1=	-129	
	data_f2=	789	;
#8000	data_f1=	-821	
	data_f2=	229	;
#8000	data_f1=	-1011	
	data_f2=	-424	;
#8000	data_f1=	-581	
	data_f2=	-903	;
#8000	data_f1=	204	
	data_f2=	-1010	;
#8000	data_f1=	864	
	data_f2=	-701	;
#8000	data_f1=	994	
	data_f2=	-103	;
#8000	data_f1=	515	
	data_f2=	538	;
#8000	data_f1=	-280	
	data_f2=	857	;
#8000	data_f1=	-904	
	data_f2=	981	;
#8000	data_f1=	-974	
	data_f2=	602	;
#8000	data_f1=	-448	
	data_f2=	-26	;
#8000	data_f1=	352	
	data_f2=	-643	;
#8000	data_f1=	937	
	data_f2=	-995	;
#8000	data_f1=	947	
	data_f2=	-937	;
#8000	data_f1=	376	
	data_f2=	-493	;
#8000	data_f1=	-425	
	data_f2=	153	;
#8000	data_f1=	-966	
	data_f2=	737	;
#8000	data_f1=	-916	
	data_f2=	1017	;
#8000	data_f1=	-305	
	data_f2=	878	;
#8000	data_f1=	493	
	data_f2=	376	;
#8000	data_f1=	988	
	data_f2=	-279	;
#8000	data_f1=	878	
	data_f2=	-820	;
#8000	data_f1=	229	
	data_f2=	-1023	;
#8000	data_f1=	-560	
	data_f2=	-805	;
#8000	data_f1=	-1006	
	data_f2=	-254	;
#8000	data_f1=	-836	
	data_f2=	401	;
#8000	data_f1=	-154	
	data_f2=	891	;
#8000	data_f1=	622	
	data_f2=	1014	;
#8000	data_f1=	1017	
	data_f2=	719	;
#8000	data_f1=	789	
	data_f2=	128	;
#8000	data_f1=	77	
	data_f2=	-515	;
#8000	data_f1=	-682	
	data_f2=	-947	;
#8000	data_f1=	-1024	
	data_f2=	-988	;
#8000	data_f1=	-738	
	data_f2=	-622	;
#8000	data_f1=	-1	
	data_f2=	0	;
*/

 endmodule
