module sin_data(
	input clk,reset,
	input [11:0] select,
	output [11:0] data_sin
);

reg [11:0] data_sin_f1;
reg [11:0] data_sin_f2;

chiatan
#(
	.heso(50),
	.size(6)
)
clock_1m(
	.clk(clk),
	.reset(reset),
	.clk_out(clk_sample)
);

reg [9:0] cnt;
reg [12:0] temp;
reg tick;

always @(posedge clk or negedge reset) begin
	if(~reset) begin
		temp <= 0;
		tick <= 1'b0;
	end
	else begin
		if(temp == 4999) begin
			tick <= 1'b1;
			temp <= temp + 1'b1;
		end
		else begin
			temp <= temp + 1'b1;
		end
	end
end

always @(posedge clk_sample or negedge reset) begin
	if(~reset) begin
		cnt <= 0;
	end
	else if(cnt == 999) begin
		cnt <= 0;
	end
	else if(tick)begin
		cnt <= cnt + 1'b1;
	end
	else begin
		cnt <= cnt;
	end
end

always @(*) begin
	if(tick) begin
		case(cnt)
		0	:	data_sin_f1 = 	2253	;
		1	:	data_sin_f1 = 	2456	;
		2	:	data_sin_f1 = 	2656	;
		3	:	data_sin_f1 = 	2849	;
		4	:	data_sin_f1 = 	3034	;
		5	:	data_sin_f1 = 	3209	;
		6	:	data_sin_f1 = 	3372	;
		7	:	data_sin_f1 = 	3522	;
		8	:	data_sin_f1 = 	3657	;
		9	:	data_sin_f1 = 	3776	;
		10	:	data_sin_f1 = 	3878	;
		11	:	data_sin_f1 = 	3961	;
		12	:	data_sin_f1 = 	4024	;
		13	:	data_sin_f1 = 	4068	;
		14	:	data_sin_f1 = 	4091	;
		15	:	data_sin_f1 = 	4094	;
		16	:	data_sin_f1 = 	4075	;
		17	:	data_sin_f1 = 	4037	;
		18	:	data_sin_f1 = 	3978	;
		19	:	data_sin_f1 = 	3900	;
		20	:	data_sin_f1 = 	3803	;
		21	:	data_sin_f1 = 	3689	;
		22	:	data_sin_f1 = 	3558	;
		23	:	data_sin_f1 = 	3411	;
		24	:	data_sin_f1 = 	3251	;
		25	:	data_sin_f1 = 	3079	;
		26	:	data_sin_f1 = 	2896	;
		27	:	data_sin_f1 = 	2705	;
		28	:	data_sin_f1 = 	2507	;
		29	:	data_sin_f1 = 	2304	;
		30	:	data_sin_f1 = 	2099	;
		31	:	data_sin_f1 = 	1893	;
		32	:	data_sin_f1 = 	1689	;
		33	:	data_sin_f1 = 	1489	;
		34	:	data_sin_f1 = 	1294	;
		35	:	data_sin_f1 = 	1107	;
		36	:	data_sin_f1 = 	929	;
		37	:	data_sin_f1 = 	762	;
		38	:	data_sin_f1 = 	609	;
		39	:	data_sin_f1 = 	470	;
		40	:	data_sin_f1 = 	347	;
		41	:	data_sin_f1 = 	241	;
		42	:	data_sin_f1 = 	153	;
		43	:	data_sin_f1 = 	85	;
		44	:	data_sin_f1 = 	36	;
		45	:	data_sin_f1 = 	8	;
		46	:	data_sin_f1 = 	0	;
		47	:	data_sin_f1 = 	13	;
		48	:	data_sin_f1 = 	47	;
		49	:	data_sin_f1 = 	100	;
		50	:	data_sin_f1 = 	174	;
		51	:	data_sin_f1 = 	266	;
		52	:	data_sin_f1 = 	376	;
		53	:	data_sin_f1 = 	503	;
		54	:	data_sin_f1 = 	646	;
		55	:	data_sin_f1 = 	803	;
		56	:	data_sin_f1 = 	972	;
		57	:	data_sin_f1 = 	1153	;
		58	:	data_sin_f1 = 	1342	;
		59	:	data_sin_f1 = 	1538	;
		60	:	data_sin_f1 = 	1740	;
		61	:	data_sin_f1 = 	1945	;
		62	:	data_sin_f1 = 	2150	;
		63	:	data_sin_f1 = 	2355	;
		64	:	data_sin_f1 = 	2557	;
		65	:	data_sin_f1 = 	2753	;
		66	:	data_sin_f1 = 	2942	;
		67	:	data_sin_f1 = 	3123	;
		68	:	data_sin_f1 = 	3292	;
		69	:	data_sin_f1 = 	3449	;
		70	:	data_sin_f1 = 	3592	;
		71	:	data_sin_f1 = 	3719	;
		72	:	data_sin_f1 = 	3829	;
		73	:	data_sin_f1 = 	3921	;
		74	:	data_sin_f1 = 	3995	;
		75	:	data_sin_f1 = 	4048	;
		76	:	data_sin_f1 = 	4082	;
		77	:	data_sin_f1 = 	4095	;
		78	:	data_sin_f1 = 	4087	;
		79	:	data_sin_f1 = 	4059	;
		80	:	data_sin_f1 = 	4010	;
		81	:	data_sin_f1 = 	3942	;
		82	:	data_sin_f1 = 	3854	;
		83	:	data_sin_f1 = 	3748	;
		84	:	data_sin_f1 = 	3625	;
		85	:	data_sin_f1 = 	3486	;
		86	:	data_sin_f1 = 	3333	;
		87	:	data_sin_f1 = 	3166	;
		88	:	data_sin_f1 = 	2988	;
		89	:	data_sin_f1 = 	2801	;
		90	:	data_sin_f1 = 	2606	;
		91	:	data_sin_f1 = 	2406	;
		92	:	data_sin_f1 = 	2202	;
		93	:	data_sin_f1 = 	1996	;
		94	:	data_sin_f1 = 	1791	;
		95	:	data_sin_f1 = 	1588	;
		96	:	data_sin_f1 = 	1390	;
		97	:	data_sin_f1 = 	1199	;
		98	:	data_sin_f1 = 	1016	;
		99	:	data_sin_f1 = 	844	;
		100	:	data_sin_f1 = 	684	;
		101	:	data_sin_f1 = 	537	;
		102	:	data_sin_f1 = 	406	;
		103	:	data_sin_f1 = 	292	;
		104	:	data_sin_f1 = 	195	;
		105	:	data_sin_f1 = 	117	;
		106	:	data_sin_f1 = 	58	;
		107	:	data_sin_f1 = 	20	;
		108	:	data_sin_f1 = 	1	;
		109	:	data_sin_f1 = 	4	;
		110	:	data_sin_f1 = 	27	;
		111	:	data_sin_f1 = 	71	;
		112	:	data_sin_f1 = 	134	;
		113	:	data_sin_f1 = 	217	;
		114	:	data_sin_f1 = 	319	;
		115	:	data_sin_f1 = 	438	;
		116	:	data_sin_f1 = 	573	;
		117	:	data_sin_f1 = 	723	;
		118	:	data_sin_f1 = 	886	;
		119	:	data_sin_f1 = 	1061	;
		120	:	data_sin_f1 = 	1246	;
		121	:	data_sin_f1 = 	1439	;
		122	:	data_sin_f1 = 	1639	;
		123	:	data_sin_f1 = 	1842	;
		124	:	data_sin_f1 = 	2048	;
		125	:	data_sin_f1 = 	2253	;
		126	:	data_sin_f1 = 	2456	;
		127	:	data_sin_f1 = 	2656	;
		128	:	data_sin_f1 = 	2849	;
		129	:	data_sin_f1 = 	3034	;
		130	:	data_sin_f1 = 	3209	;
		131	:	data_sin_f1 = 	3372	;
		132	:	data_sin_f1 = 	3522	;
		133	:	data_sin_f1 = 	3657	;
		134	:	data_sin_f1 = 	3776	;
		135	:	data_sin_f1 = 	3878	;
		136	:	data_sin_f1 = 	3961	;
		137	:	data_sin_f1 = 	4024	;
		138	:	data_sin_f1 = 	4068	;
		139	:	data_sin_f1 = 	4091	;
		140	:	data_sin_f1 = 	4094	;
		141	:	data_sin_f1 = 	4075	;
		142	:	data_sin_f1 = 	4037	;
		143	:	data_sin_f1 = 	3978	;
		144	:	data_sin_f1 = 	3900	;
		145	:	data_sin_f1 = 	3803	;
		146	:	data_sin_f1 = 	3689	;
		147	:	data_sin_f1 = 	3558	;
		148	:	data_sin_f1 = 	3411	;
		149	:	data_sin_f1 = 	3251	;
		150	:	data_sin_f1 = 	3079	;
		151	:	data_sin_f1 = 	2896	;
		152	:	data_sin_f1 = 	2705	;
		153	:	data_sin_f1 = 	2507	;
		154	:	data_sin_f1 = 	2304	;
		155	:	data_sin_f1 = 	2099	;
		156	:	data_sin_f1 = 	1893	;
		157	:	data_sin_f1 = 	1689	;
		158	:	data_sin_f1 = 	1489	;
		159	:	data_sin_f1 = 	1294	;
		160	:	data_sin_f1 = 	1107	;
		161	:	data_sin_f1 = 	929	;
		162	:	data_sin_f1 = 	762	;
		163	:	data_sin_f1 = 	609	;
		164	:	data_sin_f1 = 	470	;
		165	:	data_sin_f1 = 	347	;
		166	:	data_sin_f1 = 	241	;
		167	:	data_sin_f1 = 	153	;
		168	:	data_sin_f1 = 	85	;
		169	:	data_sin_f1 = 	36	;
		170	:	data_sin_f1 = 	8	;
		171	:	data_sin_f1 = 	0	;
		172	:	data_sin_f1 = 	13	;
		173	:	data_sin_f1 = 	47	;
		174	:	data_sin_f1 = 	100	;
		175	:	data_sin_f1 = 	174	;
		176	:	data_sin_f1 = 	266	;
		177	:	data_sin_f1 = 	376	;
		178	:	data_sin_f1 = 	503	;
		179	:	data_sin_f1 = 	646	;
		180	:	data_sin_f1 = 	803	;
		181	:	data_sin_f1 = 	972	;
		182	:	data_sin_f1 = 	1153	;
		183	:	data_sin_f1 = 	1342	;
		184	:	data_sin_f1 = 	1538	;
		185	:	data_sin_f1 = 	1740	;
		186	:	data_sin_f1 = 	1945	;
		187	:	data_sin_f1 = 	2150	;
		188	:	data_sin_f1 = 	2355	;
		189	:	data_sin_f1 = 	2557	;
		190	:	data_sin_f1 = 	2753	;
		191	:	data_sin_f1 = 	2942	;
		192	:	data_sin_f1 = 	3123	;
		193	:	data_sin_f1 = 	3292	;
		194	:	data_sin_f1 = 	3449	;
		195	:	data_sin_f1 = 	3592	;
		196	:	data_sin_f1 = 	3719	;
		197	:	data_sin_f1 = 	3829	;
		198	:	data_sin_f1 = 	3921	;
		199	:	data_sin_f1 = 	3995	;
		200	:	data_sin_f1 = 	4048	;
		201	:	data_sin_f1 = 	4082	;
		202	:	data_sin_f1 = 	4095	;
		203	:	data_sin_f1 = 	4087	;
		204	:	data_sin_f1 = 	4059	;
		205	:	data_sin_f1 = 	4010	;
		206	:	data_sin_f1 = 	3942	;
		207	:	data_sin_f1 = 	3854	;
		208	:	data_sin_f1 = 	3748	;
		209	:	data_sin_f1 = 	3625	;
		210	:	data_sin_f1 = 	3486	;
		211	:	data_sin_f1 = 	3333	;
		212	:	data_sin_f1 = 	3166	;
		213	:	data_sin_f1 = 	2988	;
		214	:	data_sin_f1 = 	2801	;
		215	:	data_sin_f1 = 	2606	;
		216	:	data_sin_f1 = 	2406	;
		217	:	data_sin_f1 = 	2202	;
		218	:	data_sin_f1 = 	1996	;
		219	:	data_sin_f1 = 	1791	;
		220	:	data_sin_f1 = 	1588	;
		221	:	data_sin_f1 = 	1390	;
		222	:	data_sin_f1 = 	1199	;
		223	:	data_sin_f1 = 	1016	;
		224	:	data_sin_f1 = 	844	;
		225	:	data_sin_f1 = 	684	;
		226	:	data_sin_f1 = 	537	;
		227	:	data_sin_f1 = 	406	;
		228	:	data_sin_f1 = 	292	;
		229	:	data_sin_f1 = 	195	;
		230	:	data_sin_f1 = 	117	;
		231	:	data_sin_f1 = 	58	;
		232	:	data_sin_f1 = 	20	;
		233	:	data_sin_f1 = 	1	;
		234	:	data_sin_f1 = 	4	;
		235	:	data_sin_f1 = 	27	;
		236	:	data_sin_f1 = 	71	;
		237	:	data_sin_f1 = 	134	;
		238	:	data_sin_f1 = 	217	;
		239	:	data_sin_f1 = 	319	;
		240	:	data_sin_f1 = 	438	;
		241	:	data_sin_f1 = 	573	;
		242	:	data_sin_f1 = 	723	;
		243	:	data_sin_f1 = 	886	;
		244	:	data_sin_f1 = 	1061	;
		245	:	data_sin_f1 = 	1246	;
		246	:	data_sin_f1 = 	1439	;
		247	:	data_sin_f1 = 	1639	;
		248	:	data_sin_f1 = 	1842	;
		249	:	data_sin_f1 = 	2048	;
		250	:	data_sin_f1 = 	2253	;
		251	:	data_sin_f1 = 	2456	;
		252	:	data_sin_f1 = 	2656	;
		253	:	data_sin_f1 = 	2849	;
		254	:	data_sin_f1 = 	3034	;
		255	:	data_sin_f1 = 	3209	;
		256	:	data_sin_f1 = 	3372	;
		257	:	data_sin_f1 = 	3522	;
		258	:	data_sin_f1 = 	3657	;
		259	:	data_sin_f1 = 	3776	;
		260	:	data_sin_f1 = 	3878	;
		261	:	data_sin_f1 = 	3961	;
		262	:	data_sin_f1 = 	4024	;
		263	:	data_sin_f1 = 	4068	;
		264	:	data_sin_f1 = 	4091	;
		265	:	data_sin_f1 = 	4094	;
		266	:	data_sin_f1 = 	4075	;
		267	:	data_sin_f1 = 	4037	;
		268	:	data_sin_f1 = 	3978	;
		269	:	data_sin_f1 = 	3900	;
		270	:	data_sin_f1 = 	3803	;
		271	:	data_sin_f1 = 	3689	;
		272	:	data_sin_f1 = 	3558	;
		273	:	data_sin_f1 = 	3411	;
		274	:	data_sin_f1 = 	3251	;
		275	:	data_sin_f1 = 	3079	;
		276	:	data_sin_f1 = 	2896	;
		277	:	data_sin_f1 = 	2705	;
		278	:	data_sin_f1 = 	2507	;
		279	:	data_sin_f1 = 	2304	;
		280	:	data_sin_f1 = 	2099	;
		281	:	data_sin_f1 = 	1893	;
		282	:	data_sin_f1 = 	1689	;
		283	:	data_sin_f1 = 	1489	;
		284	:	data_sin_f1 = 	1294	;
		285	:	data_sin_f1 = 	1107	;
		286	:	data_sin_f1 = 	929	;
		287	:	data_sin_f1 = 	762	;
		288	:	data_sin_f1 = 	609	;
		289	:	data_sin_f1 = 	470	;
		290	:	data_sin_f1 = 	347	;
		291	:	data_sin_f1 = 	241	;
		292	:	data_sin_f1 = 	153	;
		293	:	data_sin_f1 = 	85	;
		294	:	data_sin_f1 = 	36	;
		295	:	data_sin_f1 = 	8	;
		296	:	data_sin_f1 = 	0	;
		297	:	data_sin_f1 = 	13	;
		298	:	data_sin_f1 = 	47	;
		299	:	data_sin_f1 = 	100	;
		300	:	data_sin_f1 = 	174	;
		301	:	data_sin_f1 = 	266	;
		302	:	data_sin_f1 = 	376	;
		303	:	data_sin_f1 = 	503	;
		304	:	data_sin_f1 = 	646	;
		305	:	data_sin_f1 = 	803	;
		306	:	data_sin_f1 = 	972	;
		307	:	data_sin_f1 = 	1153	;
		308	:	data_sin_f1 = 	1342	;
		309	:	data_sin_f1 = 	1538	;
		310	:	data_sin_f1 = 	1740	;
		311	:	data_sin_f1 = 	1945	;
		312	:	data_sin_f1 = 	2150	;
		313	:	data_sin_f1 = 	2355	;
		314	:	data_sin_f1 = 	2557	;
		315	:	data_sin_f1 = 	2753	;
		316	:	data_sin_f1 = 	2942	;
		317	:	data_sin_f1 = 	3123	;
		318	:	data_sin_f1 = 	3292	;
		319	:	data_sin_f1 = 	3449	;
		320	:	data_sin_f1 = 	3592	;
		321	:	data_sin_f1 = 	3719	;
		322	:	data_sin_f1 = 	3829	;
		323	:	data_sin_f1 = 	3921	;
		324	:	data_sin_f1 = 	3995	;
		325	:	data_sin_f1 = 	4048	;
		326	:	data_sin_f1 = 	4082	;
		327	:	data_sin_f1 = 	4095	;
		328	:	data_sin_f1 = 	4087	;
		329	:	data_sin_f1 = 	4059	;
		330	:	data_sin_f1 = 	4010	;
		331	:	data_sin_f1 = 	3942	;
		332	:	data_sin_f1 = 	3854	;
		333	:	data_sin_f1 = 	3748	;
		334	:	data_sin_f1 = 	3625	;
		335	:	data_sin_f1 = 	3486	;
		336	:	data_sin_f1 = 	3333	;
		337	:	data_sin_f1 = 	3166	;
		338	:	data_sin_f1 = 	2988	;
		339	:	data_sin_f1 = 	2801	;
		340	:	data_sin_f1 = 	2606	;
		341	:	data_sin_f1 = 	2406	;
		342	:	data_sin_f1 = 	2202	;
		343	:	data_sin_f1 = 	1996	;
		344	:	data_sin_f1 = 	1791	;
		345	:	data_sin_f1 = 	1588	;
		346	:	data_sin_f1 = 	1390	;
		347	:	data_sin_f1 = 	1199	;
		348	:	data_sin_f1 = 	1016	;
		349	:	data_sin_f1 = 	844	;
		350	:	data_sin_f1 = 	684	;
		351	:	data_sin_f1 = 	537	;
		352	:	data_sin_f1 = 	406	;
		353	:	data_sin_f1 = 	292	;
		354	:	data_sin_f1 = 	195	;
		355	:	data_sin_f1 = 	117	;
		356	:	data_sin_f1 = 	58	;
		357	:	data_sin_f1 = 	20	;
		358	:	data_sin_f1 = 	1	;
		359	:	data_sin_f1 = 	4	;
		360	:	data_sin_f1 = 	27	;
		361	:	data_sin_f1 = 	71	;
		362	:	data_sin_f1 = 	134	;
		363	:	data_sin_f1 = 	217	;
		364	:	data_sin_f1 = 	319	;
		365	:	data_sin_f1 = 	438	;
		366	:	data_sin_f1 = 	573	;
		367	:	data_sin_f1 = 	723	;
		368	:	data_sin_f1 = 	886	;
		369	:	data_sin_f1 = 	1061	;
		370	:	data_sin_f1 = 	1246	;
		371	:	data_sin_f1 = 	1439	;
		372	:	data_sin_f1 = 	1639	;
		373	:	data_sin_f1 = 	1842	;
		374	:	data_sin_f1 = 	2048	;
		375	:	data_sin_f1 = 	2253	;
		376	:	data_sin_f1 = 	2456	;
		377	:	data_sin_f1 = 	2656	;
		378	:	data_sin_f1 = 	2849	;
		379	:	data_sin_f1 = 	3034	;
		380	:	data_sin_f1 = 	3209	;
		381	:	data_sin_f1 = 	3372	;
		382	:	data_sin_f1 = 	3522	;
		383	:	data_sin_f1 = 	3657	;
		384	:	data_sin_f1 = 	3776	;
		385	:	data_sin_f1 = 	3878	;
		386	:	data_sin_f1 = 	3961	;
		387	:	data_sin_f1 = 	4024	;
		388	:	data_sin_f1 = 	4068	;
		389	:	data_sin_f1 = 	4091	;
		390	:	data_sin_f1 = 	4094	;
		391	:	data_sin_f1 = 	4075	;
		392	:	data_sin_f1 = 	4037	;
		393	:	data_sin_f1 = 	3978	;
		394	:	data_sin_f1 = 	3900	;
		395	:	data_sin_f1 = 	3803	;
		396	:	data_sin_f1 = 	3689	;
		397	:	data_sin_f1 = 	3558	;
		398	:	data_sin_f1 = 	3411	;
		399	:	data_sin_f1 = 	3251	;
		400	:	data_sin_f1 = 	3079	;
		401	:	data_sin_f1 = 	2896	;
		402	:	data_sin_f1 = 	2705	;
		403	:	data_sin_f1 = 	2507	;
		404	:	data_sin_f1 = 	2304	;
		405	:	data_sin_f1 = 	2099	;
		406	:	data_sin_f1 = 	1893	;
		407	:	data_sin_f1 = 	1689	;
		408	:	data_sin_f1 = 	1489	;
		409	:	data_sin_f1 = 	1294	;
		410	:	data_sin_f1 = 	1107	;
		411	:	data_sin_f1 = 	929	;
		412	:	data_sin_f1 = 	762	;
		413	:	data_sin_f1 = 	609	;
		414	:	data_sin_f1 = 	470	;
		415	:	data_sin_f1 = 	347	;
		416	:	data_sin_f1 = 	241	;
		417	:	data_sin_f1 = 	153	;
		418	:	data_sin_f1 = 	85	;
		419	:	data_sin_f1 = 	36	;
		420	:	data_sin_f1 = 	8	;
		421	:	data_sin_f1 = 	0	;
		422	:	data_sin_f1 = 	13	;
		423	:	data_sin_f1 = 	47	;
		424	:	data_sin_f1 = 	100	;
		425	:	data_sin_f1 = 	174	;
		426	:	data_sin_f1 = 	266	;
		427	:	data_sin_f1 = 	376	;
		428	:	data_sin_f1 = 	503	;
		429	:	data_sin_f1 = 	646	;
		430	:	data_sin_f1 = 	803	;
		431	:	data_sin_f1 = 	972	;
		432	:	data_sin_f1 = 	1153	;
		433	:	data_sin_f1 = 	1342	;
		434	:	data_sin_f1 = 	1538	;
		435	:	data_sin_f1 = 	1740	;
		436	:	data_sin_f1 = 	1945	;
		437	:	data_sin_f1 = 	2150	;
		438	:	data_sin_f1 = 	2355	;
		439	:	data_sin_f1 = 	2557	;
		440	:	data_sin_f1 = 	2753	;
		441	:	data_sin_f1 = 	2942	;
		442	:	data_sin_f1 = 	3123	;
		443	:	data_sin_f1 = 	3292	;
		444	:	data_sin_f1 = 	3449	;
		445	:	data_sin_f1 = 	3592	;
		446	:	data_sin_f1 = 	3719	;
		447	:	data_sin_f1 = 	3829	;
		448	:	data_sin_f1 = 	3921	;
		449	:	data_sin_f1 = 	3995	;
		450	:	data_sin_f1 = 	4048	;
		451	:	data_sin_f1 = 	4082	;
		452	:	data_sin_f1 = 	4095	;
		453	:	data_sin_f1 = 	4087	;
		454	:	data_sin_f1 = 	4059	;
		455	:	data_sin_f1 = 	4010	;
		456	:	data_sin_f1 = 	3942	;
		457	:	data_sin_f1 = 	3854	;
		458	:	data_sin_f1 = 	3748	;
		459	:	data_sin_f1 = 	3625	;
		460	:	data_sin_f1 = 	3486	;
		461	:	data_sin_f1 = 	3333	;
		462	:	data_sin_f1 = 	3166	;
		463	:	data_sin_f1 = 	2988	;
		464	:	data_sin_f1 = 	2801	;
		465	:	data_sin_f1 = 	2606	;
		466	:	data_sin_f1 = 	2406	;
		467	:	data_sin_f1 = 	2202	;
		468	:	data_sin_f1 = 	1996	;
		469	:	data_sin_f1 = 	1791	;
		470	:	data_sin_f1 = 	1588	;
		471	:	data_sin_f1 = 	1390	;
		472	:	data_sin_f1 = 	1199	;
		473	:	data_sin_f1 = 	1016	;
		474	:	data_sin_f1 = 	844	;
		475	:	data_sin_f1 = 	684	;
		476	:	data_sin_f1 = 	537	;
		477	:	data_sin_f1 = 	406	;
		478	:	data_sin_f1 = 	292	;
		479	:	data_sin_f1 = 	195	;
		480	:	data_sin_f1 = 	117	;
		481	:	data_sin_f1 = 	58	;
		482	:	data_sin_f1 = 	20	;
		483	:	data_sin_f1 = 	1	;
		484	:	data_sin_f1 = 	4	;
		485	:	data_sin_f1 = 	27	;
		486	:	data_sin_f1 = 	71	;
		487	:	data_sin_f1 = 	134	;
		488	:	data_sin_f1 = 	217	;
		489	:	data_sin_f1 = 	319	;
		490	:	data_sin_f1 = 	438	;
		491	:	data_sin_f1 = 	573	;
		492	:	data_sin_f1 = 	723	;
		493	:	data_sin_f1 = 	886	;
		494	:	data_sin_f1 = 	1061	;
		495	:	data_sin_f1 = 	1246	;
		496	:	data_sin_f1 = 	1439	;
		497	:	data_sin_f1 = 	1639	;
		498	:	data_sin_f1 = 	1842	;
		499	:	data_sin_f1 = 	2048	;
		500	:	data_sin_f1 = 	2253	;
		501	:	data_sin_f1 = 	2456	;
		502	:	data_sin_f1 = 	2656	;
		503	:	data_sin_f1 = 	2849	;
		504	:	data_sin_f1 = 	3034	;
		505	:	data_sin_f1 = 	3209	;
		506	:	data_sin_f1 = 	3372	;
		507	:	data_sin_f1 = 	3522	;
		508	:	data_sin_f1 = 	3657	;
		509	:	data_sin_f1 = 	3776	;
		510	:	data_sin_f1 = 	3878	;
		511	:	data_sin_f1 = 	3961	;
		512	:	data_sin_f1 = 	4024	;
		513	:	data_sin_f1 = 	4068	;
		514	:	data_sin_f1 = 	4091	;
		515	:	data_sin_f1 = 	4094	;
		516	:	data_sin_f1 = 	4075	;
		517	:	data_sin_f1 = 	4037	;
		518	:	data_sin_f1 = 	3978	;
		519	:	data_sin_f1 = 	3900	;
		520	:	data_sin_f1 = 	3803	;
		521	:	data_sin_f1 = 	3689	;
		522	:	data_sin_f1 = 	3558	;
		523	:	data_sin_f1 = 	3411	;
		524	:	data_sin_f1 = 	3251	;
		525	:	data_sin_f1 = 	3079	;
		526	:	data_sin_f1 = 	2896	;
		527	:	data_sin_f1 = 	2705	;
		528	:	data_sin_f1 = 	2507	;
		529	:	data_sin_f1 = 	2304	;
		530	:	data_sin_f1 = 	2099	;
		531	:	data_sin_f1 = 	1893	;
		532	:	data_sin_f1 = 	1689	;
		533	:	data_sin_f1 = 	1489	;
		534	:	data_sin_f1 = 	1294	;
		535	:	data_sin_f1 = 	1107	;
		536	:	data_sin_f1 = 	929	;
		537	:	data_sin_f1 = 	762	;
		538	:	data_sin_f1 = 	609	;
		539	:	data_sin_f1 = 	470	;
		540	:	data_sin_f1 = 	347	;
		541	:	data_sin_f1 = 	241	;
		542	:	data_sin_f1 = 	153	;
		543	:	data_sin_f1 = 	85	;
		544	:	data_sin_f1 = 	36	;
		545	:	data_sin_f1 = 	8	;
		546	:	data_sin_f1 = 	0	;
		547	:	data_sin_f1 = 	13	;
		548	:	data_sin_f1 = 	47	;
		549	:	data_sin_f1 = 	100	;
		550	:	data_sin_f1 = 	174	;
		551	:	data_sin_f1 = 	266	;
		552	:	data_sin_f1 = 	376	;
		553	:	data_sin_f1 = 	503	;
		554	:	data_sin_f1 = 	646	;
		555	:	data_sin_f1 = 	803	;
		556	:	data_sin_f1 = 	972	;
		557	:	data_sin_f1 = 	1153	;
		558	:	data_sin_f1 = 	1342	;
		559	:	data_sin_f1 = 	1538	;
		560	:	data_sin_f1 = 	1740	;
		561	:	data_sin_f1 = 	1945	;
		562	:	data_sin_f1 = 	2150	;
		563	:	data_sin_f1 = 	2355	;
		564	:	data_sin_f1 = 	2557	;
		565	:	data_sin_f1 = 	2753	;
		566	:	data_sin_f1 = 	2942	;
		567	:	data_sin_f1 = 	3123	;
		568	:	data_sin_f1 = 	3292	;
		569	:	data_sin_f1 = 	3449	;
		570	:	data_sin_f1 = 	3592	;
		571	:	data_sin_f1 = 	3719	;
		572	:	data_sin_f1 = 	3829	;
		573	:	data_sin_f1 = 	3921	;
		574	:	data_sin_f1 = 	3995	;
		575	:	data_sin_f1 = 	4048	;
		576	:	data_sin_f1 = 	4082	;
		577	:	data_sin_f1 = 	4095	;
		578	:	data_sin_f1 = 	4087	;
		579	:	data_sin_f1 = 	4059	;
		580	:	data_sin_f1 = 	4010	;
		581	:	data_sin_f1 = 	3942	;
		582	:	data_sin_f1 = 	3854	;
		583	:	data_sin_f1 = 	3748	;
		584	:	data_sin_f1 = 	3625	;
		585	:	data_sin_f1 = 	3486	;
		586	:	data_sin_f1 = 	3333	;
		587	:	data_sin_f1 = 	3166	;
		588	:	data_sin_f1 = 	2988	;
		589	:	data_sin_f1 = 	2801	;
		590	:	data_sin_f1 = 	2606	;
		591	:	data_sin_f1 = 	2406	;
		592	:	data_sin_f1 = 	2202	;
		593	:	data_sin_f1 = 	1996	;
		594	:	data_sin_f1 = 	1791	;
		595	:	data_sin_f1 = 	1588	;
		596	:	data_sin_f1 = 	1390	;
		597	:	data_sin_f1 = 	1199	;
		598	:	data_sin_f1 = 	1016	;
		599	:	data_sin_f1 = 	844	;
		600	:	data_sin_f1 = 	684	;
		601	:	data_sin_f1 = 	537	;
		602	:	data_sin_f1 = 	406	;
		603	:	data_sin_f1 = 	292	;
		604	:	data_sin_f1 = 	195	;
		605	:	data_sin_f1 = 	117	;
		606	:	data_sin_f1 = 	58	;
		607	:	data_sin_f1 = 	20	;
		608	:	data_sin_f1 = 	1	;
		609	:	data_sin_f1 = 	4	;
		610	:	data_sin_f1 = 	27	;
		611	:	data_sin_f1 = 	71	;
		612	:	data_sin_f1 = 	134	;
		613	:	data_sin_f1 = 	217	;
		614	:	data_sin_f1 = 	319	;
		615	:	data_sin_f1 = 	438	;
		616	:	data_sin_f1 = 	573	;
		617	:	data_sin_f1 = 	723	;
		618	:	data_sin_f1 = 	886	;
		619	:	data_sin_f1 = 	1061	;
		620	:	data_sin_f1 = 	1246	;
		621	:	data_sin_f1 = 	1439	;
		622	:	data_sin_f1 = 	1639	;
		623	:	data_sin_f1 = 	1842	;
		624	:	data_sin_f1 = 	2048	;
		625	:	data_sin_f1 = 	2253	;
		626	:	data_sin_f1 = 	2456	;
		627	:	data_sin_f1 = 	2656	;
		628	:	data_sin_f1 = 	2849	;
		629	:	data_sin_f1 = 	3034	;
		630	:	data_sin_f1 = 	3209	;
		631	:	data_sin_f1 = 	3372	;
		632	:	data_sin_f1 = 	3522	;
		633	:	data_sin_f1 = 	3657	;
		634	:	data_sin_f1 = 	3776	;
		635	:	data_sin_f1 = 	3878	;
		636	:	data_sin_f1 = 	3961	;
		637	:	data_sin_f1 = 	4024	;
		638	:	data_sin_f1 = 	4068	;
		639	:	data_sin_f1 = 	4091	;
		640	:	data_sin_f1 = 	4094	;
		641	:	data_sin_f1 = 	4075	;
		642	:	data_sin_f1 = 	4037	;
		643	:	data_sin_f1 = 	3978	;
		644	:	data_sin_f1 = 	3900	;
		645	:	data_sin_f1 = 	3803	;
		646	:	data_sin_f1 = 	3689	;
		647	:	data_sin_f1 = 	3558	;
		648	:	data_sin_f1 = 	3411	;
		649	:	data_sin_f1 = 	3251	;
		650	:	data_sin_f1 = 	3079	;
		651	:	data_sin_f1 = 	2896	;
		652	:	data_sin_f1 = 	2705	;
		653	:	data_sin_f1 = 	2507	;
		654	:	data_sin_f1 = 	2304	;
		655	:	data_sin_f1 = 	2099	;
		656	:	data_sin_f1 = 	1893	;
		657	:	data_sin_f1 = 	1689	;
		658	:	data_sin_f1 = 	1489	;
		659	:	data_sin_f1 = 	1294	;
		660	:	data_sin_f1 = 	1107	;
		661	:	data_sin_f1 = 	929	;
		662	:	data_sin_f1 = 	762	;
		663	:	data_sin_f1 = 	609	;
		664	:	data_sin_f1 = 	470	;
		665	:	data_sin_f1 = 	347	;
		666	:	data_sin_f1 = 	241	;
		667	:	data_sin_f1 = 	153	;
		668	:	data_sin_f1 = 	85	;
		669	:	data_sin_f1 = 	36	;
		670	:	data_sin_f1 = 	8	;
		671	:	data_sin_f1 = 	0	;
		672	:	data_sin_f1 = 	13	;
		673	:	data_sin_f1 = 	47	;
		674	:	data_sin_f1 = 	100	;
		675	:	data_sin_f1 = 	174	;
		676	:	data_sin_f1 = 	266	;
		677	:	data_sin_f1 = 	376	;
		678	:	data_sin_f1 = 	503	;
		679	:	data_sin_f1 = 	646	;
		680	:	data_sin_f1 = 	803	;
		681	:	data_sin_f1 = 	972	;
		682	:	data_sin_f1 = 	1153	;
		683	:	data_sin_f1 = 	1342	;
		684	:	data_sin_f1 = 	1538	;
		685	:	data_sin_f1 = 	1740	;
		686	:	data_sin_f1 = 	1945	;
		687	:	data_sin_f1 = 	2150	;
		688	:	data_sin_f1 = 	2355	;
		689	:	data_sin_f1 = 	2557	;
		690	:	data_sin_f1 = 	2753	;
		691	:	data_sin_f1 = 	2942	;
		692	:	data_sin_f1 = 	3123	;
		693	:	data_sin_f1 = 	3292	;
		694	:	data_sin_f1 = 	3449	;
		695	:	data_sin_f1 = 	3592	;
		696	:	data_sin_f1 = 	3719	;
		697	:	data_sin_f1 = 	3829	;
		698	:	data_sin_f1 = 	3921	;
		699	:	data_sin_f1 = 	3995	;
		700	:	data_sin_f1 = 	4048	;
		701	:	data_sin_f1 = 	4082	;
		702	:	data_sin_f1 = 	4095	;
		703	:	data_sin_f1 = 	4087	;
		704	:	data_sin_f1 = 	4059	;
		705	:	data_sin_f1 = 	4010	;
		706	:	data_sin_f1 = 	3942	;
		707	:	data_sin_f1 = 	3854	;
		708	:	data_sin_f1 = 	3748	;
		709	:	data_sin_f1 = 	3625	;
		710	:	data_sin_f1 = 	3486	;
		711	:	data_sin_f1 = 	3333	;
		712	:	data_sin_f1 = 	3166	;
		713	:	data_sin_f1 = 	2988	;
		714	:	data_sin_f1 = 	2801	;
		715	:	data_sin_f1 = 	2606	;
		716	:	data_sin_f1 = 	2406	;
		717	:	data_sin_f1 = 	2202	;
		718	:	data_sin_f1 = 	1996	;
		719	:	data_sin_f1 = 	1791	;
		720	:	data_sin_f1 = 	1588	;
		721	:	data_sin_f1 = 	1390	;
		722	:	data_sin_f1 = 	1199	;
		723	:	data_sin_f1 = 	1016	;
		724	:	data_sin_f1 = 	844	;
		725	:	data_sin_f1 = 	684	;
		726	:	data_sin_f1 = 	537	;
		727	:	data_sin_f1 = 	406	;
		728	:	data_sin_f1 = 	292	;
		729	:	data_sin_f1 = 	195	;
		730	:	data_sin_f1 = 	117	;
		731	:	data_sin_f1 = 	58	;
		732	:	data_sin_f1 = 	20	;
		733	:	data_sin_f1 = 	1	;
		734	:	data_sin_f1 = 	4	;
		735	:	data_sin_f1 = 	27	;
		736	:	data_sin_f1 = 	71	;
		737	:	data_sin_f1 = 	134	;
		738	:	data_sin_f1 = 	217	;
		739	:	data_sin_f1 = 	319	;
		740	:	data_sin_f1 = 	438	;
		741	:	data_sin_f1 = 	573	;
		742	:	data_sin_f1 = 	723	;
		743	:	data_sin_f1 = 	886	;
		744	:	data_sin_f1 = 	1061	;
		745	:	data_sin_f1 = 	1246	;
		746	:	data_sin_f1 = 	1439	;
		747	:	data_sin_f1 = 	1639	;
		748	:	data_sin_f1 = 	1842	;
		749	:	data_sin_f1 = 	2047	;
		750	:	data_sin_f1 = 	2253	;
		751	:	data_sin_f1 = 	2456	;
		752	:	data_sin_f1 = 	2656	;
		753	:	data_sin_f1 = 	2849	;
		754	:	data_sin_f1 = 	3034	;
		755	:	data_sin_f1 = 	3209	;
		756	:	data_sin_f1 = 	3372	;
		757	:	data_sin_f1 = 	3522	;
		758	:	data_sin_f1 = 	3657	;
		759	:	data_sin_f1 = 	3776	;
		760	:	data_sin_f1 = 	3878	;
		761	:	data_sin_f1 = 	3961	;
		762	:	data_sin_f1 = 	4024	;
		763	:	data_sin_f1 = 	4068	;
		764	:	data_sin_f1 = 	4091	;
		765	:	data_sin_f1 = 	4094	;
		766	:	data_sin_f1 = 	4075	;
		767	:	data_sin_f1 = 	4037	;
		768	:	data_sin_f1 = 	3978	;
		769	:	data_sin_f1 = 	3900	;
		770	:	data_sin_f1 = 	3803	;
		771	:	data_sin_f1 = 	3689	;
		772	:	data_sin_f1 = 	3558	;
		773	:	data_sin_f1 = 	3411	;
		774	:	data_sin_f1 = 	3251	;
		775	:	data_sin_f1 = 	3079	;
		776	:	data_sin_f1 = 	2896	;
		777	:	data_sin_f1 = 	2705	;
		778	:	data_sin_f1 = 	2507	;
		779	:	data_sin_f1 = 	2304	;
		780	:	data_sin_f1 = 	2099	;
		781	:	data_sin_f1 = 	1893	;
		782	:	data_sin_f1 = 	1689	;
		783	:	data_sin_f1 = 	1489	;
		784	:	data_sin_f1 = 	1294	;
		785	:	data_sin_f1 = 	1107	;
		786	:	data_sin_f1 = 	929	;
		787	:	data_sin_f1 = 	762	;
		788	:	data_sin_f1 = 	609	;
		789	:	data_sin_f1 = 	470	;
		790	:	data_sin_f1 = 	347	;
		791	:	data_sin_f1 = 	241	;
		792	:	data_sin_f1 = 	153	;
		793	:	data_sin_f1 = 	85	;
		794	:	data_sin_f1 = 	36	;
		795	:	data_sin_f1 = 	8	;
		796	:	data_sin_f1 = 	0	;
		797	:	data_sin_f1 = 	13	;
		798	:	data_sin_f1 = 	47	;
		799	:	data_sin_f1 = 	100	;
		800	:	data_sin_f1 = 	174	;
		801	:	data_sin_f1 = 	266	;
		802	:	data_sin_f1 = 	376	;
		803	:	data_sin_f1 = 	503	;
		804	:	data_sin_f1 = 	646	;
		805	:	data_sin_f1 = 	803	;
		806	:	data_sin_f1 = 	972	;
		807	:	data_sin_f1 = 	1153	;
		808	:	data_sin_f1 = 	1342	;
		809	:	data_sin_f1 = 	1538	;
		810	:	data_sin_f1 = 	1740	;
		811	:	data_sin_f1 = 	1945	;
		812	:	data_sin_f1 = 	2150	;
		813	:	data_sin_f1 = 	2355	;
		814	:	data_sin_f1 = 	2557	;
		815	:	data_sin_f1 = 	2753	;
		816	:	data_sin_f1 = 	2942	;
		817	:	data_sin_f1 = 	3123	;
		818	:	data_sin_f1 = 	3292	;
		819	:	data_sin_f1 = 	3449	;
		820	:	data_sin_f1 = 	3592	;
		821	:	data_sin_f1 = 	3719	;
		822	:	data_sin_f1 = 	3829	;
		823	:	data_sin_f1 = 	3921	;
		824	:	data_sin_f1 = 	3995	;
		825	:	data_sin_f1 = 	4048	;
		826	:	data_sin_f1 = 	4082	;
		827	:	data_sin_f1 = 	4095	;
		828	:	data_sin_f1 = 	4087	;
		829	:	data_sin_f1 = 	4059	;
		830	:	data_sin_f1 = 	4010	;
		831	:	data_sin_f1 = 	3942	;
		832	:	data_sin_f1 = 	3854	;
		833	:	data_sin_f1 = 	3748	;
		834	:	data_sin_f1 = 	3625	;
		835	:	data_sin_f1 = 	3486	;
		836	:	data_sin_f1 = 	3333	;
		837	:	data_sin_f1 = 	3166	;
		838	:	data_sin_f1 = 	2988	;
		839	:	data_sin_f1 = 	2801	;
		840	:	data_sin_f1 = 	2606	;
		841	:	data_sin_f1 = 	2406	;
		842	:	data_sin_f1 = 	2202	;
		843	:	data_sin_f1 = 	1996	;
		844	:	data_sin_f1 = 	1791	;
		845	:	data_sin_f1 = 	1588	;
		846	:	data_sin_f1 = 	1390	;
		847	:	data_sin_f1 = 	1199	;
		848	:	data_sin_f1 = 	1016	;
		849	:	data_sin_f1 = 	844	;
		850	:	data_sin_f1 = 	684	;
		851	:	data_sin_f1 = 	537	;
		852	:	data_sin_f1 = 	406	;
		853	:	data_sin_f1 = 	292	;
		854	:	data_sin_f1 = 	195	;
		855	:	data_sin_f1 = 	117	;
		856	:	data_sin_f1 = 	58	;
		857	:	data_sin_f1 = 	20	;
		858	:	data_sin_f1 = 	1	;
		859	:	data_sin_f1 = 	4	;
		860	:	data_sin_f1 = 	27	;
		861	:	data_sin_f1 = 	71	;
		862	:	data_sin_f1 = 	134	;
		863	:	data_sin_f1 = 	217	;
		864	:	data_sin_f1 = 	319	;
		865	:	data_sin_f1 = 	438	;
		866	:	data_sin_f1 = 	573	;
		867	:	data_sin_f1 = 	723	;
		868	:	data_sin_f1 = 	886	;
		869	:	data_sin_f1 = 	1061	;
		870	:	data_sin_f1 = 	1246	;
		871	:	data_sin_f1 = 	1439	;
		872	:	data_sin_f1 = 	1639	;
		873	:	data_sin_f1 = 	1842	;
		874	:	data_sin_f1 = 	2047	;
		875	:	data_sin_f1 = 	2253	;
		876	:	data_sin_f1 = 	2456	;
		877	:	data_sin_f1 = 	2656	;
		878	:	data_sin_f1 = 	2849	;
		879	:	data_sin_f1 = 	3034	;
		880	:	data_sin_f1 = 	3209	;
		881	:	data_sin_f1 = 	3372	;
		882	:	data_sin_f1 = 	3522	;
		883	:	data_sin_f1 = 	3657	;
		884	:	data_sin_f1 = 	3776	;
		885	:	data_sin_f1 = 	3878	;
		886	:	data_sin_f1 = 	3961	;
		887	:	data_sin_f1 = 	4024	;
		888	:	data_sin_f1 = 	4068	;
		889	:	data_sin_f1 = 	4091	;
		890	:	data_sin_f1 = 	4094	;
		891	:	data_sin_f1 = 	4075	;
		892	:	data_sin_f1 = 	4037	;
		893	:	data_sin_f1 = 	3978	;
		894	:	data_sin_f1 = 	3900	;
		895	:	data_sin_f1 = 	3803	;
		896	:	data_sin_f1 = 	3689	;
		897	:	data_sin_f1 = 	3558	;
		898	:	data_sin_f1 = 	3411	;
		899	:	data_sin_f1 = 	3251	;
		900	:	data_sin_f1 = 	3079	;
		901	:	data_sin_f1 = 	2896	;
		902	:	data_sin_f1 = 	2705	;
		903	:	data_sin_f1 = 	2507	;
		904	:	data_sin_f1 = 	2304	;
		905	:	data_sin_f1 = 	2099	;
		906	:	data_sin_f1 = 	1893	;
		907	:	data_sin_f1 = 	1689	;
		908	:	data_sin_f1 = 	1489	;
		909	:	data_sin_f1 = 	1294	;
		910	:	data_sin_f1 = 	1107	;
		911	:	data_sin_f1 = 	929	;
		912	:	data_sin_f1 = 	762	;
		913	:	data_sin_f1 = 	609	;
		914	:	data_sin_f1 = 	470	;
		915	:	data_sin_f1 = 	347	;
		916	:	data_sin_f1 = 	241	;
		917	:	data_sin_f1 = 	153	;
		918	:	data_sin_f1 = 	85	;
		919	:	data_sin_f1 = 	36	;
		920	:	data_sin_f1 = 	8	;
		921	:	data_sin_f1 = 	0	;
		922	:	data_sin_f1 = 	13	;
		923	:	data_sin_f1 = 	47	;
		924	:	data_sin_f1 = 	100	;
		925	:	data_sin_f1 = 	174	;
		926	:	data_sin_f1 = 	266	;
		927	:	data_sin_f1 = 	376	;
		928	:	data_sin_f1 = 	503	;
		929	:	data_sin_f1 = 	646	;
		930	:	data_sin_f1 = 	803	;
		931	:	data_sin_f1 = 	972	;
		932	:	data_sin_f1 = 	1153	;
		933	:	data_sin_f1 = 	1342	;
		934	:	data_sin_f1 = 	1538	;
		935	:	data_sin_f1 = 	1740	;
		936	:	data_sin_f1 = 	1945	;
		937	:	data_sin_f1 = 	2150	;
		938	:	data_sin_f1 = 	2355	;
		939	:	data_sin_f1 = 	2557	;
		940	:	data_sin_f1 = 	2753	;
		941	:	data_sin_f1 = 	2942	;
		942	:	data_sin_f1 = 	3123	;
		943	:	data_sin_f1 = 	3292	;
		944	:	data_sin_f1 = 	3449	;
		945	:	data_sin_f1 = 	3592	;
		946	:	data_sin_f1 = 	3719	;
		947	:	data_sin_f1 = 	3829	;
		948	:	data_sin_f1 = 	3921	;
		949	:	data_sin_f1 = 	3995	;
		950	:	data_sin_f1 = 	4048	;
		951	:	data_sin_f1 = 	4082	;
		952	:	data_sin_f1 = 	4095	;
		953	:	data_sin_f1 = 	4087	;
		954	:	data_sin_f1 = 	4059	;
		955	:	data_sin_f1 = 	4010	;
		956	:	data_sin_f1 = 	3942	;
		957	:	data_sin_f1 = 	3854	;
		958	:	data_sin_f1 = 	3748	;
		959	:	data_sin_f1 = 	3625	;
		960	:	data_sin_f1 = 	3486	;
		961	:	data_sin_f1 = 	3333	;
		962	:	data_sin_f1 = 	3166	;
		963	:	data_sin_f1 = 	2988	;
		964	:	data_sin_f1 = 	2801	;
		965	:	data_sin_f1 = 	2606	;
		966	:	data_sin_f1 = 	2406	;
		967	:	data_sin_f1 = 	2202	;
		968	:	data_sin_f1 = 	1996	;
		969	:	data_sin_f1 = 	1791	;
		970	:	data_sin_f1 = 	1588	;
		971	:	data_sin_f1 = 	1390	;
		972	:	data_sin_f1 = 	1199	;
		973	:	data_sin_f1 = 	1016	;
		974	:	data_sin_f1 = 	844	;
		975	:	data_sin_f1 = 	684	;
		976	:	data_sin_f1 = 	537	;
		977	:	data_sin_f1 = 	406	;
		978	:	data_sin_f1 = 	292	;
		979	:	data_sin_f1 = 	195	;
		980	:	data_sin_f1 = 	117	;
		981	:	data_sin_f1 = 	58	;
		982	:	data_sin_f1 = 	20	;
		983	:	data_sin_f1 = 	1	;
		984	:	data_sin_f1 = 	4	;
		985	:	data_sin_f1 = 	27	;
		986	:	data_sin_f1 = 	71	;
		987	:	data_sin_f1 = 	134	;
		988	:	data_sin_f1 = 	217	;
		989	:	data_sin_f1 = 	319	;
		990	:	data_sin_f1 = 	438	;
		991	:	data_sin_f1 = 	573	;
		992	:	data_sin_f1 = 	723	;
		993	:	data_sin_f1 = 	886	;
		994	:	data_sin_f1 = 	1061	;
		995	:	data_sin_f1 = 	1246	;
		996	:	data_sin_f1 = 	1439	;
		997	:	data_sin_f1 = 	1639	;
		998	:	data_sin_f1 = 	1842	;
		999	:	data_sin_f1 = 	2047	;
		default: data_sin_f1 = 2047;
	endcase
	end
	else
		data_sin_f1 = 2047;
end

always @(*) begin
	if(tick) begin
		case(cnt)
		0	:	data_sin_f2 = 	2215	;
1	:	data_sin_f2 = 	2380	;
2	:	data_sin_f2 = 	2544	;
3	:	data_sin_f2 = 	2705	;
4	:	data_sin_f2 = 	2861	;
5	:	data_sin_f2 = 	3011	;
6	:	data_sin_f2 = 	3155	;
7	:	data_sin_f2 = 	3292	;
8	:	data_sin_f2 = 	3421	;
9	:	data_sin_f2 = 	3540	;
10	:	data_sin_f2 = 	3649	;
11	:	data_sin_f2 = 	3748	;
12	:	data_sin_f2 = 	3836	;
13	:	data_sin_f2 = 	3911	;
14	:	data_sin_f2 = 	3974	;
15	:	data_sin_f2 = 	4024	;
16	:	data_sin_f2 = 	4061	;
17	:	data_sin_f2 = 	4085	;
18	:	data_sin_f2 = 	4095	;
19	:	data_sin_f2 = 	4091	;
20	:	data_sin_f2 = 	4074	;
21	:	data_sin_f2 = 	4043	;
22	:	data_sin_f2 = 	3999	;
23	:	data_sin_f2 = 	3942	;
24	:	data_sin_f2 = 	3872	;
25	:	data_sin_f2 = 	3790	;
26	:	data_sin_f2 = 	3696	;
27	:	data_sin_f2 = 	3592	;
28	:	data_sin_f2 = 	3477	;
29	:	data_sin_f2 = 	3353	;
30	:	data_sin_f2 = 	3220	;
31	:	data_sin_f2 = 	3079	;
32	:	data_sin_f2 = 	2931	;
33	:	data_sin_f2 = 	2777	;
34	:	data_sin_f2 = 	2619	;
35	:	data_sin_f2 = 	2456	;
36	:	data_sin_f2 = 	2291	;
37	:	data_sin_f2 = 	2125	;
38	:	data_sin_f2 = 	1957	;
39	:	data_sin_f2 = 	1791	;
40	:	data_sin_f2 = 	1626	;
41	:	data_sin_f2 = 	1464	;
42	:	data_sin_f2 = 	1306	;
43	:	data_sin_f2 = 	1153	;
44	:	data_sin_f2 = 	1005	;
45	:	data_sin_f2 = 	865	;
46	:	data_sin_f2 = 	732	;
47	:	data_sin_f2 = 	609	;
48	:	data_sin_f2 = 	495	;
49	:	data_sin_f2 = 	391	;
50	:	data_sin_f2 = 	298	;
51	:	data_sin_f2 = 	217	;
52	:	data_sin_f2 = 	149	;
53	:	data_sin_f2 = 	92	;
54	:	data_sin_f2 = 	49	;
55	:	data_sin_f2 = 	20	;
56	:	data_sin_f2 = 	3	;
57	:	data_sin_f2 = 	1	;
58	:	data_sin_f2 = 	12	;
59	:	data_sin_f2 = 	36	;
60	:	data_sin_f2 = 	74	;
61	:	data_sin_f2 = 	125	;
62	:	data_sin_f2 = 	189	;
63	:	data_sin_f2 = 	266	;
64	:	data_sin_f2 = 	354	;
65	:	data_sin_f2 = 	454	;
66	:	data_sin_f2 = 	564	;
67	:	data_sin_f2 = 	684	;
68	:	data_sin_f2 = 	813	;
69	:	data_sin_f2 = 	950	;
70	:	data_sin_f2 = 	1095	;
71	:	data_sin_f2 = 	1246	;
72	:	data_sin_f2 = 	1403	;
73	:	data_sin_f2 = 	1563	;
74	:	data_sin_f2 = 	1727	;
75	:	data_sin_f2 = 	1893	;
76	:	data_sin_f2 = 	2060	;
77	:	data_sin_f2 = 	2227	;
78	:	data_sin_f2 = 	2393	;
79	:	data_sin_f2 = 	2557	;
80	:	data_sin_f2 = 	2717	;
81	:	data_sin_f2 = 	2872	;
82	:	data_sin_f2 = 	3023	;
83	:	data_sin_f2 = 	3166	;
84	:	data_sin_f2 = 	3302	;
85	:	data_sin_f2 = 	3430	;
86	:	data_sin_f2 = 	3549	;
87	:	data_sin_f2 = 	3657	;
88	:	data_sin_f2 = 	3755	;
89	:	data_sin_f2 = 	3842	;
90	:	data_sin_f2 = 	3916	;
91	:	data_sin_f2 = 	3978	;
92	:	data_sin_f2 = 	4027	;
93	:	data_sin_f2 = 	4063	;
94	:	data_sin_f2 = 	4086	;
95	:	data_sin_f2 = 	4095	;
96	:	data_sin_f2 = 	4090	;
97	:	data_sin_f2 = 	4072	;
98	:	data_sin_f2 = 	4040	;
99	:	data_sin_f2 = 	3995	;
100	:	data_sin_f2 = 	3937	;
101	:	data_sin_f2 = 	3866	;
102	:	data_sin_f2 = 	3783	;
103	:	data_sin_f2 = 	3689	;
104	:	data_sin_f2 = 	3583	;
105	:	data_sin_f2 = 	3468	;
106	:	data_sin_f2 = 	3343	;
107	:	data_sin_f2 = 	3209	;
108	:	data_sin_f2 = 	3068	;
109	:	data_sin_f2 = 	2919	;
110	:	data_sin_f2 = 	2765	;
111	:	data_sin_f2 = 	2606	;
112	:	data_sin_f2 = 	2444	;
113	:	data_sin_f2 = 	2279	;
114	:	data_sin_f2 = 	2112	;
115	:	data_sin_f2 = 	1945	;
116	:	data_sin_f2 = 	1778	;
117	:	data_sin_f2 = 	1613	;
118	:	data_sin_f2 = 	1452	;
119	:	data_sin_f2 = 	1294	;
120	:	data_sin_f2 = 	1141	;
121	:	data_sin_f2 = 	994	;
122	:	data_sin_f2 = 	854	;
123	:	data_sin_f2 = 	723	;
124	:	data_sin_f2 = 	600	;
125	:	data_sin_f2 = 	486	;
126	:	data_sin_f2 = 	384	;
127	:	data_sin_f2 = 	292	;
128	:	data_sin_f2 = 	212	;
129	:	data_sin_f2 = 	144	;
130	:	data_sin_f2 = 	89	;
131	:	data_sin_f2 = 	47	;
132	:	data_sin_f2 = 	18	;
133	:	data_sin_f2 = 	3	;
134	:	data_sin_f2 = 	1	;
135	:	data_sin_f2 = 	13	;
136	:	data_sin_f2 = 	39	;
137	:	data_sin_f2 = 	78	;
138	:	data_sin_f2 = 	130	;
139	:	data_sin_f2 = 	195	;
140	:	data_sin_f2 = 	272	;
141	:	data_sin_f2 = 	361	;
142	:	data_sin_f2 = 	462	;
143	:	data_sin_f2 = 	573	;
144	:	data_sin_f2 = 	693	;
145	:	data_sin_f2 = 	823	;
146	:	data_sin_f2 = 	961	;
147	:	data_sin_f2 = 	1107	;
148	:	data_sin_f2 = 	1258	;
149	:	data_sin_f2 = 	1415	;
150	:	data_sin_f2 = 	1576	;
151	:	data_sin_f2 = 	1740	;
152	:	data_sin_f2 = 	1906	;
153	:	data_sin_f2 = 	2073	;
154	:	data_sin_f2 = 	2240	;
155	:	data_sin_f2 = 	2406	;
156	:	data_sin_f2 = 	2569	;
157	:	data_sin_f2 = 	2729	;
158	:	data_sin_f2 = 	2884	;
159	:	data_sin_f2 = 	3034	;
160	:	data_sin_f2 = 	3177	;
161	:	data_sin_f2 = 	3313	;
162	:	data_sin_f2 = 	3440	;
163	:	data_sin_f2 = 	3558	;
164	:	data_sin_f2 = 	3665	;
165	:	data_sin_f2 = 	3762	;
166	:	data_sin_f2 = 	3848	;
167	:	data_sin_f2 = 	3921	;
168	:	data_sin_f2 = 	3983	;
169	:	data_sin_f2 = 	4031	;
170	:	data_sin_f2 = 	4066	;
171	:	data_sin_f2 = 	4087	;
172	:	data_sin_f2 = 	4095	;
173	:	data_sin_f2 = 	4089	;
174	:	data_sin_f2 = 	4070	;
175	:	data_sin_f2 = 	4037	;
176	:	data_sin_f2 = 	3991	;
177	:	data_sin_f2 = 	3932	;
178	:	data_sin_f2 = 	3860	;
179	:	data_sin_f2 = 	3776	;
180	:	data_sin_f2 = 	3681	;
181	:	data_sin_f2 = 	3575	;
182	:	data_sin_f2 = 	3458	;
183	:	data_sin_f2 = 	3333	;
184	:	data_sin_f2 = 	3198	;
185	:	data_sin_f2 = 	3056	;
186	:	data_sin_f2 = 	2908	;
187	:	data_sin_f2 = 	2753	;
188	:	data_sin_f2 = 	2594	;
189	:	data_sin_f2 = 	2431	;
190	:	data_sin_f2 = 	2266	;
191	:	data_sin_f2 = 	2099	;
192	:	data_sin_f2 = 	1932	;
193	:	data_sin_f2 = 	1765	;
194	:	data_sin_f2 = 	1601	;
195	:	data_sin_f2 = 	1439	;
196	:	data_sin_f2 = 	1282	;
197	:	data_sin_f2 = 	1129	;
198	:	data_sin_f2 = 	983	;
199	:	data_sin_f2 = 	844	;
200	:	data_sin_f2 = 	713	;
201	:	data_sin_f2 = 	591	;
202	:	data_sin_f2 = 	478	;
203	:	data_sin_f2 = 	376	;
204	:	data_sin_f2 = 	285	;
205	:	data_sin_f2 = 	206	;
206	:	data_sin_f2 = 	139	;
207	:	data_sin_f2 = 	85	;
208	:	data_sin_f2 = 	44	;
209	:	data_sin_f2 = 	16	;
210	:	data_sin_f2 = 	2	;
211	:	data_sin_f2 = 	1	;
212	:	data_sin_f2 = 	15	;
213	:	data_sin_f2 = 	41	;
214	:	data_sin_f2 = 	81	;
215	:	data_sin_f2 = 	134	;
216	:	data_sin_f2 = 	200	;
217	:	data_sin_f2 = 	279	;
218	:	data_sin_f2 = 	369	;
219	:	data_sin_f2 = 	470	;
220	:	data_sin_f2 = 	582	;
221	:	data_sin_f2 = 	703	;
222	:	data_sin_f2 = 	834	;
223	:	data_sin_f2 = 	972	;
224	:	data_sin_f2 = 	1118	;
225	:	data_sin_f2 = 	1270	;
226	:	data_sin_f2 = 	1427	;
227	:	data_sin_f2 = 	1588	;
228	:	data_sin_f2 = 	1753	;
229	:	data_sin_f2 = 	1919	;
230	:	data_sin_f2 = 	2086	;
231	:	data_sin_f2 = 	2253	;
232	:	data_sin_f2 = 	2419	;
233	:	data_sin_f2 = 	2582	;
234	:	data_sin_f2 = 	2741	;
235	:	data_sin_f2 = 	2896	;
236	:	data_sin_f2 = 	3045	;
237	:	data_sin_f2 = 	3188	;
238	:	data_sin_f2 = 	3323	;
239	:	data_sin_f2 = 	3449	;
240	:	data_sin_f2 = 	3566	;
241	:	data_sin_f2 = 	3673	;
242	:	data_sin_f2 = 	3769	;
243	:	data_sin_f2 = 	3854	;
244	:	data_sin_f2 = 	3927	;
245	:	data_sin_f2 = 	3987	;
246	:	data_sin_f2 = 	4034	;
247	:	data_sin_f2 = 	4068	;
248	:	data_sin_f2 = 	4088	;
249	:	data_sin_f2 = 	4095	;
250	:	data_sin_f2 = 	4088	;
251	:	data_sin_f2 = 	4068	;
252	:	data_sin_f2 = 	4034	;
253	:	data_sin_f2 = 	3987	;
254	:	data_sin_f2 = 	3927	;
255	:	data_sin_f2 = 	3854	;
256	:	data_sin_f2 = 	3769	;
257	:	data_sin_f2 = 	3673	;
258	:	data_sin_f2 = 	3566	;
259	:	data_sin_f2 = 	3449	;
260	:	data_sin_f2 = 	3323	;
261	:	data_sin_f2 = 	3188	;
262	:	data_sin_f2 = 	3045	;
263	:	data_sin_f2 = 	2896	;
264	:	data_sin_f2 = 	2741	;
265	:	data_sin_f2 = 	2582	;
266	:	data_sin_f2 = 	2419	;
267	:	data_sin_f2 = 	2253	;
268	:	data_sin_f2 = 	2086	;
269	:	data_sin_f2 = 	1919	;
270	:	data_sin_f2 = 	1753	;
271	:	data_sin_f2 = 	1588	;
272	:	data_sin_f2 = 	1427	;
273	:	data_sin_f2 = 	1270	;
274	:	data_sin_f2 = 	1118	;
275	:	data_sin_f2 = 	972	;
276	:	data_sin_f2 = 	834	;
277	:	data_sin_f2 = 	703	;
278	:	data_sin_f2 = 	582	;
279	:	data_sin_f2 = 	470	;
280	:	data_sin_f2 = 	369	;
281	:	data_sin_f2 = 	279	;
282	:	data_sin_f2 = 	200	;
283	:	data_sin_f2 = 	134	;
284	:	data_sin_f2 = 	81	;
285	:	data_sin_f2 = 	41	;
286	:	data_sin_f2 = 	15	;
287	:	data_sin_f2 = 	1	;
288	:	data_sin_f2 = 	2	;
289	:	data_sin_f2 = 	16	;
290	:	data_sin_f2 = 	44	;
291	:	data_sin_f2 = 	85	;
292	:	data_sin_f2 = 	139	;
293	:	data_sin_f2 = 	206	;
294	:	data_sin_f2 = 	285	;
295	:	data_sin_f2 = 	376	;
296	:	data_sin_f2 = 	478	;
297	:	data_sin_f2 = 	591	;
298	:	data_sin_f2 = 	713	;
299	:	data_sin_f2 = 	844	;
300	:	data_sin_f2 = 	983	;
301	:	data_sin_f2 = 	1129	;
302	:	data_sin_f2 = 	1282	;
303	:	data_sin_f2 = 	1439	;
304	:	data_sin_f2 = 	1601	;
305	:	data_sin_f2 = 	1765	;
306	:	data_sin_f2 = 	1932	;
307	:	data_sin_f2 = 	2099	;
308	:	data_sin_f2 = 	2266	;
309	:	data_sin_f2 = 	2431	;
310	:	data_sin_f2 = 	2594	;
311	:	data_sin_f2 = 	2753	;
312	:	data_sin_f2 = 	2908	;
313	:	data_sin_f2 = 	3056	;
314	:	data_sin_f2 = 	3198	;
315	:	data_sin_f2 = 	3333	;
316	:	data_sin_f2 = 	3458	;
317	:	data_sin_f2 = 	3575	;
318	:	data_sin_f2 = 	3681	;
319	:	data_sin_f2 = 	3776	;
320	:	data_sin_f2 = 	3860	;
321	:	data_sin_f2 = 	3932	;
322	:	data_sin_f2 = 	3991	;
323	:	data_sin_f2 = 	4037	;
324	:	data_sin_f2 = 	4070	;
325	:	data_sin_f2 = 	4089	;
326	:	data_sin_f2 = 	4095	;
327	:	data_sin_f2 = 	4087	;
328	:	data_sin_f2 = 	4066	;
329	:	data_sin_f2 = 	4031	;
330	:	data_sin_f2 = 	3983	;
331	:	data_sin_f2 = 	3921	;
332	:	data_sin_f2 = 	3848	;
333	:	data_sin_f2 = 	3762	;
334	:	data_sin_f2 = 	3665	;
335	:	data_sin_f2 = 	3558	;
336	:	data_sin_f2 = 	3440	;
337	:	data_sin_f2 = 	3313	;
338	:	data_sin_f2 = 	3177	;
339	:	data_sin_f2 = 	3034	;
340	:	data_sin_f2 = 	2884	;
341	:	data_sin_f2 = 	2729	;
342	:	data_sin_f2 = 	2569	;
343	:	data_sin_f2 = 	2406	;
344	:	data_sin_f2 = 	2240	;
345	:	data_sin_f2 = 	2073	;
346	:	data_sin_f2 = 	1906	;
347	:	data_sin_f2 = 	1740	;
348	:	data_sin_f2 = 	1576	;
349	:	data_sin_f2 = 	1415	;
350	:	data_sin_f2 = 	1258	;
351	:	data_sin_f2 = 	1107	;
352	:	data_sin_f2 = 	961	;
353	:	data_sin_f2 = 	823	;
354	:	data_sin_f2 = 	693	;
355	:	data_sin_f2 = 	573	;
356	:	data_sin_f2 = 	462	;
357	:	data_sin_f2 = 	361	;
358	:	data_sin_f2 = 	272	;
359	:	data_sin_f2 = 	195	;
360	:	data_sin_f2 = 	130	;
361	:	data_sin_f2 = 	78	;
362	:	data_sin_f2 = 	39	;
363	:	data_sin_f2 = 	13	;
364	:	data_sin_f2 = 	1	;
365	:	data_sin_f2 = 	3	;
366	:	data_sin_f2 = 	18	;
367	:	data_sin_f2 = 	47	;
368	:	data_sin_f2 = 	89	;
369	:	data_sin_f2 = 	144	;
370	:	data_sin_f2 = 	212	;
371	:	data_sin_f2 = 	292	;
372	:	data_sin_f2 = 	384	;
373	:	data_sin_f2 = 	486	;
374	:	data_sin_f2 = 	600	;
375	:	data_sin_f2 = 	723	;
376	:	data_sin_f2 = 	854	;
377	:	data_sin_f2 = 	994	;
378	:	data_sin_f2 = 	1141	;
379	:	data_sin_f2 = 	1294	;
380	:	data_sin_f2 = 	1452	;
381	:	data_sin_f2 = 	1613	;
382	:	data_sin_f2 = 	1778	;
383	:	data_sin_f2 = 	1945	;
384	:	data_sin_f2 = 	2112	;
385	:	data_sin_f2 = 	2279	;
386	:	data_sin_f2 = 	2444	;
387	:	data_sin_f2 = 	2606	;
388	:	data_sin_f2 = 	2765	;
389	:	data_sin_f2 = 	2919	;
390	:	data_sin_f2 = 	3068	;
391	:	data_sin_f2 = 	3209	;
392	:	data_sin_f2 = 	3343	;
393	:	data_sin_f2 = 	3468	;
394	:	data_sin_f2 = 	3583	;
395	:	data_sin_f2 = 	3689	;
396	:	data_sin_f2 = 	3783	;
397	:	data_sin_f2 = 	3866	;
398	:	data_sin_f2 = 	3937	;
399	:	data_sin_f2 = 	3995	;
400	:	data_sin_f2 = 	4040	;
401	:	data_sin_f2 = 	4072	;
402	:	data_sin_f2 = 	4090	;
403	:	data_sin_f2 = 	4095	;
404	:	data_sin_f2 = 	4086	;
405	:	data_sin_f2 = 	4063	;
406	:	data_sin_f2 = 	4027	;
407	:	data_sin_f2 = 	3978	;
408	:	data_sin_f2 = 	3916	;
409	:	data_sin_f2 = 	3842	;
410	:	data_sin_f2 = 	3755	;
411	:	data_sin_f2 = 	3657	;
412	:	data_sin_f2 = 	3549	;
413	:	data_sin_f2 = 	3430	;
414	:	data_sin_f2 = 	3302	;
415	:	data_sin_f2 = 	3166	;
416	:	data_sin_f2 = 	3023	;
417	:	data_sin_f2 = 	2872	;
418	:	data_sin_f2 = 	2717	;
419	:	data_sin_f2 = 	2557	;
420	:	data_sin_f2 = 	2393	;
421	:	data_sin_f2 = 	2227	;
422	:	data_sin_f2 = 	2060	;
423	:	data_sin_f2 = 	1893	;
424	:	data_sin_f2 = 	1727	;
425	:	data_sin_f2 = 	1563	;
426	:	data_sin_f2 = 	1403	;
427	:	data_sin_f2 = 	1246	;
428	:	data_sin_f2 = 	1095	;
429	:	data_sin_f2 = 	950	;
430	:	data_sin_f2 = 	813	;
431	:	data_sin_f2 = 	684	;
432	:	data_sin_f2 = 	564	;
433	:	data_sin_f2 = 	454	;
434	:	data_sin_f2 = 	354	;
435	:	data_sin_f2 = 	266	;
436	:	data_sin_f2 = 	189	;
437	:	data_sin_f2 = 	125	;
438	:	data_sin_f2 = 	74	;
439	:	data_sin_f2 = 	36	;
440	:	data_sin_f2 = 	12	;
441	:	data_sin_f2 = 	1	;
442	:	data_sin_f2 = 	3	;
443	:	data_sin_f2 = 	20	;
444	:	data_sin_f2 = 	49	;
445	:	data_sin_f2 = 	92	;
446	:	data_sin_f2 = 	149	;
447	:	data_sin_f2 = 	217	;
448	:	data_sin_f2 = 	298	;
449	:	data_sin_f2 = 	391	;
450	:	data_sin_f2 = 	495	;
451	:	data_sin_f2 = 	609	;
452	:	data_sin_f2 = 	732	;
453	:	data_sin_f2 = 	865	;
454	:	data_sin_f2 = 	1005	;
455	:	data_sin_f2 = 	1153	;
456	:	data_sin_f2 = 	1306	;
457	:	data_sin_f2 = 	1464	;
458	:	data_sin_f2 = 	1626	;
459	:	data_sin_f2 = 	1791	;
460	:	data_sin_f2 = 	1957	;
461	:	data_sin_f2 = 	2125	;
462	:	data_sin_f2 = 	2291	;
463	:	data_sin_f2 = 	2456	;
464	:	data_sin_f2 = 	2619	;
465	:	data_sin_f2 = 	2777	;
466	:	data_sin_f2 = 	2931	;
467	:	data_sin_f2 = 	3079	;
468	:	data_sin_f2 = 	3220	;
469	:	data_sin_f2 = 	3353	;
470	:	data_sin_f2 = 	3477	;
471	:	data_sin_f2 = 	3592	;
472	:	data_sin_f2 = 	3696	;
473	:	data_sin_f2 = 	3790	;
474	:	data_sin_f2 = 	3872	;
475	:	data_sin_f2 = 	3942	;
476	:	data_sin_f2 = 	3999	;
477	:	data_sin_f2 = 	4043	;
478	:	data_sin_f2 = 	4074	;
479	:	data_sin_f2 = 	4091	;
480	:	data_sin_f2 = 	4095	;
481	:	data_sin_f2 = 	4085	;
482	:	data_sin_f2 = 	4061	;
483	:	data_sin_f2 = 	4024	;
484	:	data_sin_f2 = 	3974	;
485	:	data_sin_f2 = 	3911	;
486	:	data_sin_f2 = 	3836	;
487	:	data_sin_f2 = 	3748	;
488	:	data_sin_f2 = 	3649	;
489	:	data_sin_f2 = 	3540	;
490	:	data_sin_f2 = 	3421	;
491	:	data_sin_f2 = 	3292	;
492	:	data_sin_f2 = 	3155	;
493	:	data_sin_f2 = 	3011	;
494	:	data_sin_f2 = 	2861	;
495	:	data_sin_f2 = 	2705	;
496	:	data_sin_f2 = 	2544	;
497	:	data_sin_f2 = 	2380	;
498	:	data_sin_f2 = 	2215	;
499	:	data_sin_f2 = 	2048	;
500	:	data_sin_f2 = 	1880	;
501	:	data_sin_f2 = 	1715	;
502	:	data_sin_f2 = 	1551	;
503	:	data_sin_f2 = 	1390	;
504	:	data_sin_f2 = 	1234	;
505	:	data_sin_f2 = 	1084	;
506	:	data_sin_f2 = 	940	;
507	:	data_sin_f2 = 	803	;
508	:	data_sin_f2 = 	674	;
509	:	data_sin_f2 = 	555	;
510	:	data_sin_f2 = 	446	;
511	:	data_sin_f2 = 	347	;
512	:	data_sin_f2 = 	259	;
513	:	data_sin_f2 = 	184	;
514	:	data_sin_f2 = 	121	;
515	:	data_sin_f2 = 	71	;
516	:	data_sin_f2 = 	34	;
517	:	data_sin_f2 = 	10	;
518	:	data_sin_f2 = 	0	;
519	:	data_sin_f2 = 	4	;
520	:	data_sin_f2 = 	21	;
521	:	data_sin_f2 = 	52	;
522	:	data_sin_f2 = 	96	;
523	:	data_sin_f2 = 	153	;
524	:	data_sin_f2 = 	223	;
525	:	data_sin_f2 = 	305	;
526	:	data_sin_f2 = 	399	;
527	:	data_sin_f2 = 	503	;
528	:	data_sin_f2 = 	618	;
529	:	data_sin_f2 = 	742	;
530	:	data_sin_f2 = 	875	;
531	:	data_sin_f2 = 	1016	;
532	:	data_sin_f2 = 	1164	;
533	:	data_sin_f2 = 	1318	;
534	:	data_sin_f2 = 	1476	;
535	:	data_sin_f2 = 	1639	;
536	:	data_sin_f2 = 	1804	;
537	:	data_sin_f2 = 	1970	;
538	:	data_sin_f2 = 	2138	;
539	:	data_sin_f2 = 	2304	;
540	:	data_sin_f2 = 	2469	;
541	:	data_sin_f2 = 	2631	;
542	:	data_sin_f2 = 	2789	;
543	:	data_sin_f2 = 	2942	;
544	:	data_sin_f2 = 	3090	;
545	:	data_sin_f2 = 	3230	;
546	:	data_sin_f2 = 	3363	;
547	:	data_sin_f2 = 	3486	;
548	:	data_sin_f2 = 	3600	;
549	:	data_sin_f2 = 	3704	;
550	:	data_sin_f2 = 	3797	;
551	:	data_sin_f2 = 	3878	;
552	:	data_sin_f2 = 	3946	;
553	:	data_sin_f2 = 	4003	;
554	:	data_sin_f2 = 	4046	;
555	:	data_sin_f2 = 	4075	;
556	:	data_sin_f2 = 	4092	;
557	:	data_sin_f2 = 	4094	;
558	:	data_sin_f2 = 	4083	;
559	:	data_sin_f2 = 	4059	;
560	:	data_sin_f2 = 	4021	;
561	:	data_sin_f2 = 	3970	;
562	:	data_sin_f2 = 	3906	;
563	:	data_sin_f2 = 	3829	;
564	:	data_sin_f2 = 	3741	;
565	:	data_sin_f2 = 	3641	;
566	:	data_sin_f2 = 	3531	;
567	:	data_sin_f2 = 	3411	;
568	:	data_sin_f2 = 	3282	;
569	:	data_sin_f2 = 	3145	;
570	:	data_sin_f2 = 	3000	;
571	:	data_sin_f2 = 	2849	;
572	:	data_sin_f2 = 	2692	;
573	:	data_sin_f2 = 	2532	;
574	:	data_sin_f2 = 	2368	;
575	:	data_sin_f2 = 	2202	;
576	:	data_sin_f2 = 	2035	;
577	:	data_sin_f2 = 	1868	;
578	:	data_sin_f2 = 	1702	;
579	:	data_sin_f2 = 	1538	;
580	:	data_sin_f2 = 	1378	;
581	:	data_sin_f2 = 	1223	;
582	:	data_sin_f2 = 	1072	;
583	:	data_sin_f2 = 	929	;
584	:	data_sin_f2 = 	793	;
585	:	data_sin_f2 = 	665	;
586	:	data_sin_f2 = 	546	;
587	:	data_sin_f2 = 	438	;
588	:	data_sin_f2 = 	340	;
589	:	data_sin_f2 = 	253	;
590	:	data_sin_f2 = 	179	;
591	:	data_sin_f2 = 	117	;
592	:	data_sin_f2 = 	68	;
593	:	data_sin_f2 = 	32	;
594	:	data_sin_f2 = 	9	;
595	:	data_sin_f2 = 	0	;
596	:	data_sin_f2 = 	5	;
597	:	data_sin_f2 = 	23	;
598	:	data_sin_f2 = 	55	;
599	:	data_sin_f2 = 	100	;
600	:	data_sin_f2 = 	158	;
601	:	data_sin_f2 = 	229	;
602	:	data_sin_f2 = 	312	;
603	:	data_sin_f2 = 	406	;
604	:	data_sin_f2 = 	512	;
605	:	data_sin_f2 = 	627	;
606	:	data_sin_f2 = 	752	;
607	:	data_sin_f2 = 	886	;
608	:	data_sin_f2 = 	1027	;
609	:	data_sin_f2 = 	1176	;
610	:	data_sin_f2 = 	1330	;
611	:	data_sin_f2 = 	1489	;
612	:	data_sin_f2 = 	1651	;
613	:	data_sin_f2 = 	1816	;
614	:	data_sin_f2 = 	1983	;
615	:	data_sin_f2 = 	2150	;
616	:	data_sin_f2 = 	2317	;
617	:	data_sin_f2 = 	2482	;
618	:	data_sin_f2 = 	2643	;
619	:	data_sin_f2 = 	2801	;
620	:	data_sin_f2 = 	2954	;
621	:	data_sin_f2 = 	3101	;
622	:	data_sin_f2 = 	3241	;
623	:	data_sin_f2 = 	3372	;
624	:	data_sin_f2 = 	3495	;
625	:	data_sin_f2 = 	3609	;
626	:	data_sin_f2 = 	3711	;
627	:	data_sin_f2 = 	3803	;
628	:	data_sin_f2 = 	3883	;
629	:	data_sin_f2 = 	3951	;
630	:	data_sin_f2 = 	4006	;
631	:	data_sin_f2 = 	4048	;
632	:	data_sin_f2 = 	4077	;
633	:	data_sin_f2 = 	4092	;
634	:	data_sin_f2 = 	4094	;
635	:	data_sin_f2 = 	4082	;
636	:	data_sin_f2 = 	4056	;
637	:	data_sin_f2 = 	4017	;
638	:	data_sin_f2 = 	3965	;
639	:	data_sin_f2 = 	3900	;
640	:	data_sin_f2 = 	3823	;
641	:	data_sin_f2 = 	3734	;
642	:	data_sin_f2 = 	3633	;
643	:	data_sin_f2 = 	3522	;
644	:	data_sin_f2 = 	3402	;
645	:	data_sin_f2 = 	3272	;
646	:	data_sin_f2 = 	3134	;
647	:	data_sin_f2 = 	2988	;
648	:	data_sin_f2 = 	2837	;
649	:	data_sin_f2 = 	2680	;
650	:	data_sin_f2 = 	2519	;
651	:	data_sin_f2 = 	2355	;
652	:	data_sin_f2 = 	2189	;
653	:	data_sin_f2 = 	2022	;
654	:	data_sin_f2 = 	1855	;
655	:	data_sin_f2 = 	1689	;
656	:	data_sin_f2 = 	1526	;
657	:	data_sin_f2 = 	1366	;
658	:	data_sin_f2 = 	1211	;
659	:	data_sin_f2 = 	1061	;
660	:	data_sin_f2 = 	918	;
661	:	data_sin_f2 = 	782	;
662	:	data_sin_f2 = 	655	;
663	:	data_sin_f2 = 	537	;
664	:	data_sin_f2 = 	430	;
665	:	data_sin_f2 = 	333	;
666	:	data_sin_f2 = 	247	;
667	:	data_sin_f2 = 	174	;
668	:	data_sin_f2 = 	112	;
669	:	data_sin_f2 = 	64	;
670	:	data_sin_f2 = 	29	;
671	:	data_sin_f2 = 	8	;
672	:	data_sin_f2 = 	0	;
673	:	data_sin_f2 = 	6	;
674	:	data_sin_f2 = 	25	;
675	:	data_sin_f2 = 	58	;
676	:	data_sin_f2 = 	104	;
677	:	data_sin_f2 = 	163	;
678	:	data_sin_f2 = 	235	;
679	:	data_sin_f2 = 	319	;
680	:	data_sin_f2 = 	414	;
681	:	data_sin_f2 = 	520	;
682	:	data_sin_f2 = 	637	;
683	:	data_sin_f2 = 	762	;
684	:	data_sin_f2 = 	897	;
685	:	data_sin_f2 = 	1039	;
686	:	data_sin_f2 = 	1187	;
687	:	data_sin_f2 = 	1342	;
688	:	data_sin_f2 = 	1501	;
689	:	data_sin_f2 = 	1664	;
690	:	data_sin_f2 = 	1829	;
691	:	data_sin_f2 = 	1996	;
692	:	data_sin_f2 = 	2163	;
693	:	data_sin_f2 = 	2330	;
694	:	data_sin_f2 = 	2494	;
695	:	data_sin_f2 = 	2656	;
696	:	data_sin_f2 = 	2813	;
697	:	data_sin_f2 = 	2966	;
698	:	data_sin_f2 = 	3112	;
699	:	data_sin_f2 = 	3251	;
700	:	data_sin_f2 = 	3382	;
701	:	data_sin_f2 = 	3504	;
702	:	data_sin_f2 = 	3617	;
703	:	data_sin_f2 = 	3719	;
704	:	data_sin_f2 = 	3810	;
705	:	data_sin_f2 = 	3889	;
706	:	data_sin_f2 = 	3956	;
707	:	data_sin_f2 = 	4010	;
708	:	data_sin_f2 = 	4051	;
709	:	data_sin_f2 = 	4079	;
710	:	data_sin_f2 = 	4093	;
711	:	data_sin_f2 = 	4094	;
712	:	data_sin_f2 = 	4080	;
713	:	data_sin_f2 = 	4054	;
714	:	data_sin_f2 = 	4014	;
715	:	data_sin_f2 = 	3961	;
716	:	data_sin_f2 = 	3895	;
717	:	data_sin_f2 = 	3816	;
718	:	data_sin_f2 = 	3726	;
719	:	data_sin_f2 = 	3625	;
720	:	data_sin_f2 = 	3513	;
721	:	data_sin_f2 = 	3392	;
722	:	data_sin_f2 = 	3261	;
723	:	data_sin_f2 = 	3123	;
724	:	data_sin_f2 = 	2977	;
725	:	data_sin_f2 = 	2825	;
726	:	data_sin_f2 = 	2668	;
727	:	data_sin_f2 = 	2507	;
728	:	data_sin_f2 = 	2342	;
729	:	data_sin_f2 = 	2176	;
730	:	data_sin_f2 = 	2009	;
731	:	data_sin_f2 = 	1842	;
732	:	data_sin_f2 = 	1676	;
733	:	data_sin_f2 = 	1513	;
734	:	data_sin_f2 = 	1354	;
735	:	data_sin_f2 = 	1199	;
736	:	data_sin_f2 = 	1050	;
737	:	data_sin_f2 = 	907	;
738	:	data_sin_f2 = 	772	;
739	:	data_sin_f2 = 	646	;
740	:	data_sin_f2 = 	529	;
741	:	data_sin_f2 = 	422	;
742	:	data_sin_f2 = 	326	;
743	:	data_sin_f2 = 	241	;
744	:	data_sin_f2 = 	168	;
745	:	data_sin_f2 = 	108	;
746	:	data_sin_f2 = 	61	;
747	:	data_sin_f2 = 	27	;
748	:	data_sin_f2 = 	7	;
749	:	data_sin_f2 = 	0	;
750	:	data_sin_f2 = 	7	;
751	:	data_sin_f2 = 	27	;
752	:	data_sin_f2 = 	61	;
753	:	data_sin_f2 = 	108	;
754	:	data_sin_f2 = 	168	;
755	:	data_sin_f2 = 	241	;
756	:	data_sin_f2 = 	326	;
757	:	data_sin_f2 = 	422	;
758	:	data_sin_f2 = 	529	;
759	:	data_sin_f2 = 	646	;
760	:	data_sin_f2 = 	772	;
761	:	data_sin_f2 = 	907	;
762	:	data_sin_f2 = 	1050	;
763	:	data_sin_f2 = 	1199	;
764	:	data_sin_f2 = 	1354	;
765	:	data_sin_f2 = 	1513	;
766	:	data_sin_f2 = 	1676	;
767	:	data_sin_f2 = 	1842	;
768	:	data_sin_f2 = 	2009	;
769	:	data_sin_f2 = 	2176	;
770	:	data_sin_f2 = 	2342	;
771	:	data_sin_f2 = 	2507	;
772	:	data_sin_f2 = 	2668	;
773	:	data_sin_f2 = 	2825	;
774	:	data_sin_f2 = 	2977	;
775	:	data_sin_f2 = 	3123	;
776	:	data_sin_f2 = 	3261	;
777	:	data_sin_f2 = 	3392	;
778	:	data_sin_f2 = 	3513	;
779	:	data_sin_f2 = 	3625	;
780	:	data_sin_f2 = 	3726	;
781	:	data_sin_f2 = 	3816	;
782	:	data_sin_f2 = 	3895	;
783	:	data_sin_f2 = 	3961	;
784	:	data_sin_f2 = 	4014	;
785	:	data_sin_f2 = 	4054	;
786	:	data_sin_f2 = 	4080	;
787	:	data_sin_f2 = 	4094	;
788	:	data_sin_f2 = 	4093	;
789	:	data_sin_f2 = 	4079	;
790	:	data_sin_f2 = 	4051	;
791	:	data_sin_f2 = 	4010	;
792	:	data_sin_f2 = 	3956	;
793	:	data_sin_f2 = 	3889	;
794	:	data_sin_f2 = 	3810	;
795	:	data_sin_f2 = 	3719	;
796	:	data_sin_f2 = 	3617	;
797	:	data_sin_f2 = 	3504	;
798	:	data_sin_f2 = 	3382	;
799	:	data_sin_f2 = 	3251	;
800	:	data_sin_f2 = 	3112	;
801	:	data_sin_f2 = 	2966	;
802	:	data_sin_f2 = 	2813	;
803	:	data_sin_f2 = 	2656	;
804	:	data_sin_f2 = 	2494	;
805	:	data_sin_f2 = 	2330	;
806	:	data_sin_f2 = 	2163	;
807	:	data_sin_f2 = 	1996	;
808	:	data_sin_f2 = 	1829	;
809	:	data_sin_f2 = 	1664	;
810	:	data_sin_f2 = 	1501	;
811	:	data_sin_f2 = 	1342	;
812	:	data_sin_f2 = 	1187	;
813	:	data_sin_f2 = 	1039	;
814	:	data_sin_f2 = 	897	;
815	:	data_sin_f2 = 	762	;
816	:	data_sin_f2 = 	637	;
817	:	data_sin_f2 = 	520	;
818	:	data_sin_f2 = 	414	;
819	:	data_sin_f2 = 	319	;
820	:	data_sin_f2 = 	235	;
821	:	data_sin_f2 = 	163	;
822	:	data_sin_f2 = 	104	;
823	:	data_sin_f2 = 	58	;
824	:	data_sin_f2 = 	25	;
825	:	data_sin_f2 = 	6	;
826	:	data_sin_f2 = 	0	;
827	:	data_sin_f2 = 	8	;
828	:	data_sin_f2 = 	29	;
829	:	data_sin_f2 = 	64	;
830	:	data_sin_f2 = 	112	;
831	:	data_sin_f2 = 	174	;
832	:	data_sin_f2 = 	247	;
833	:	data_sin_f2 = 	333	;
834	:	data_sin_f2 = 	430	;
835	:	data_sin_f2 = 	537	;
836	:	data_sin_f2 = 	655	;
837	:	data_sin_f2 = 	782	;
838	:	data_sin_f2 = 	918	;
839	:	data_sin_f2 = 	1061	;
840	:	data_sin_f2 = 	1211	;
841	:	data_sin_f2 = 	1366	;
842	:	data_sin_f2 = 	1526	;
843	:	data_sin_f2 = 	1689	;
844	:	data_sin_f2 = 	1855	;
845	:	data_sin_f2 = 	2022	;
846	:	data_sin_f2 = 	2189	;
847	:	data_sin_f2 = 	2355	;
848	:	data_sin_f2 = 	2519	;
849	:	data_sin_f2 = 	2680	;
850	:	data_sin_f2 = 	2837	;
851	:	data_sin_f2 = 	2988	;
852	:	data_sin_f2 = 	3134	;
853	:	data_sin_f2 = 	3272	;
854	:	data_sin_f2 = 	3402	;
855	:	data_sin_f2 = 	3522	;
856	:	data_sin_f2 = 	3633	;
857	:	data_sin_f2 = 	3734	;
858	:	data_sin_f2 = 	3823	;
859	:	data_sin_f2 = 	3900	;
860	:	data_sin_f2 = 	3965	;
861	:	data_sin_f2 = 	4017	;
862	:	data_sin_f2 = 	4056	;
863	:	data_sin_f2 = 	4082	;
864	:	data_sin_f2 = 	4094	;
865	:	data_sin_f2 = 	4092	;
866	:	data_sin_f2 = 	4077	;
867	:	data_sin_f2 = 	4048	;
868	:	data_sin_f2 = 	4006	;
869	:	data_sin_f2 = 	3951	;
870	:	data_sin_f2 = 	3883	;
871	:	data_sin_f2 = 	3803	;
872	:	data_sin_f2 = 	3711	;
873	:	data_sin_f2 = 	3609	;
874	:	data_sin_f2 = 	3495	;
875	:	data_sin_f2 = 	3372	;
876	:	data_sin_f2 = 	3241	;
877	:	data_sin_f2 = 	3101	;
878	:	data_sin_f2 = 	2954	;
879	:	data_sin_f2 = 	2801	;
880	:	data_sin_f2 = 	2643	;
881	:	data_sin_f2 = 	2482	;
882	:	data_sin_f2 = 	2317	;
883	:	data_sin_f2 = 	2150	;
884	:	data_sin_f2 = 	1983	;
885	:	data_sin_f2 = 	1816	;
886	:	data_sin_f2 = 	1651	;
887	:	data_sin_f2 = 	1489	;
888	:	data_sin_f2 = 	1330	;
889	:	data_sin_f2 = 	1176	;
890	:	data_sin_f2 = 	1027	;
891	:	data_sin_f2 = 	886	;
892	:	data_sin_f2 = 	752	;
893	:	data_sin_f2 = 	627	;
894	:	data_sin_f2 = 	512	;
895	:	data_sin_f2 = 	406	;
896	:	data_sin_f2 = 	312	;
897	:	data_sin_f2 = 	229	;
898	:	data_sin_f2 = 	158	;
899	:	data_sin_f2 = 	100	;
900	:	data_sin_f2 = 	55	;
901	:	data_sin_f2 = 	23	;
902	:	data_sin_f2 = 	5	;
903	:	data_sin_f2 = 	0	;
904	:	data_sin_f2 = 	9	;
905	:	data_sin_f2 = 	32	;
906	:	data_sin_f2 = 	68	;
907	:	data_sin_f2 = 	117	;
908	:	data_sin_f2 = 	179	;
909	:	data_sin_f2 = 	253	;
910	:	data_sin_f2 = 	340	;
911	:	data_sin_f2 = 	438	;
912	:	data_sin_f2 = 	546	;
913	:	data_sin_f2 = 	665	;
914	:	data_sin_f2 = 	793	;
915	:	data_sin_f2 = 	929	;
916	:	data_sin_f2 = 	1072	;
917	:	data_sin_f2 = 	1223	;
918	:	data_sin_f2 = 	1378	;
919	:	data_sin_f2 = 	1538	;
920	:	data_sin_f2 = 	1702	;
921	:	data_sin_f2 = 	1868	;
922	:	data_sin_f2 = 	2035	;
923	:	data_sin_f2 = 	2202	;
924	:	data_sin_f2 = 	2368	;
925	:	data_sin_f2 = 	2532	;
926	:	data_sin_f2 = 	2692	;
927	:	data_sin_f2 = 	2849	;
928	:	data_sin_f2 = 	3000	;
929	:	data_sin_f2 = 	3145	;
930	:	data_sin_f2 = 	3282	;
931	:	data_sin_f2 = 	3411	;
932	:	data_sin_f2 = 	3531	;
933	:	data_sin_f2 = 	3641	;
934	:	data_sin_f2 = 	3741	;
935	:	data_sin_f2 = 	3829	;
936	:	data_sin_f2 = 	3906	;
937	:	data_sin_f2 = 	3970	;
938	:	data_sin_f2 = 	4021	;
939	:	data_sin_f2 = 	4059	;
940	:	data_sin_f2 = 	4083	;
941	:	data_sin_f2 = 	4094	;
942	:	data_sin_f2 = 	4092	;
943	:	data_sin_f2 = 	4075	;
944	:	data_sin_f2 = 	4046	;
945	:	data_sin_f2 = 	4003	;
946	:	data_sin_f2 = 	3946	;
947	:	data_sin_f2 = 	3878	;
948	:	data_sin_f2 = 	3797	;
949	:	data_sin_f2 = 	3704	;
950	:	data_sin_f2 = 	3600	;
951	:	data_sin_f2 = 	3486	;
952	:	data_sin_f2 = 	3363	;
953	:	data_sin_f2 = 	3230	;
954	:	data_sin_f2 = 	3090	;
955	:	data_sin_f2 = 	2942	;
956	:	data_sin_f2 = 	2789	;
957	:	data_sin_f2 = 	2631	;
958	:	data_sin_f2 = 	2469	;
959	:	data_sin_f2 = 	2304	;
960	:	data_sin_f2 = 	2138	;
961	:	data_sin_f2 = 	1970	;
962	:	data_sin_f2 = 	1804	;
963	:	data_sin_f2 = 	1639	;
964	:	data_sin_f2 = 	1476	;
965	:	data_sin_f2 = 	1318	;
966	:	data_sin_f2 = 	1164	;
967	:	data_sin_f2 = 	1016	;
968	:	data_sin_f2 = 	875	;
969	:	data_sin_f2 = 	742	;
970	:	data_sin_f2 = 	618	;
971	:	data_sin_f2 = 	503	;
972	:	data_sin_f2 = 	399	;
973	:	data_sin_f2 = 	305	;
974	:	data_sin_f2 = 	223	;
975	:	data_sin_f2 = 	153	;
976	:	data_sin_f2 = 	96	;
977	:	data_sin_f2 = 	52	;
978	:	data_sin_f2 = 	21	;
979	:	data_sin_f2 = 	4	;
980	:	data_sin_f2 = 	0	;
981	:	data_sin_f2 = 	10	;
982	:	data_sin_f2 = 	34	;
983	:	data_sin_f2 = 	71	;
984	:	data_sin_f2 = 	121	;
985	:	data_sin_f2 = 	184	;
986	:	data_sin_f2 = 	259	;
987	:	data_sin_f2 = 	347	;
988	:	data_sin_f2 = 	446	;
989	:	data_sin_f2 = 	555	;
990	:	data_sin_f2 = 	674	;
991	:	data_sin_f2 = 	803	;
992	:	data_sin_f2 = 	940	;
993	:	data_sin_f2 = 	1084	;
994	:	data_sin_f2 = 	1234	;
995	:	data_sin_f2 = 	1390	;
996	:	data_sin_f2 = 	1551	;
997	:	data_sin_f2 = 	1715	;
998	:	data_sin_f2 = 	1880	;
999	:	data_sin_f2 = 	2048	;
default: data_sin_f2 = 2047;
		endcase
	end
	else begin
		data_sin_f2 = 2047;
	end
end
assign data_sin = (data_sin_f1 & select) | (data_sin_f2 & ~select);
endmodule